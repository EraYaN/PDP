---------------------------------------------------------------------
-- TITLE: Random Access Memory for Xilinx
-- AUTHOR: Steve Rhoads (rhoadss@yahoo.com)
-- DATE CREATED: 11/06/05
-- FILENAME: boot_ram.vhd
-- PROJECT: Plasma CPU core
-- COPYRIGHT: Software placed into the public domain by the author.
--    Software 'as is' without warranty.  Author liable for nothing.
-- DESCRIPTION:
--    Implements Plasma internal RAM as RAMB for Spartan 3x 
--    
--    Compile the MIPS C and assembly code into "test.axf".
--    Run convert.exe to change "test.axf" to "code.txt" which
--    will contain the hex values of the opcodes.
--    Next run "ram_image ram_xilinx.vhd code.txt ram_image.vhd",
--    to create the "ram_image.vhd" file that will have the opcodes
--    correctly placed inside the INIT_00 => strings.
--    Then include ram_image.vhd in the simulation/synthesis.
--
--    Warning:  Addresses 0x1000 - 0x1FFF are reserved for the cache
--    if the DDR cache is enabled.
---------------------------------------------------------------------
-- UPDATED: 09/07/10 Olivier Rinaudo (orinaudo@gmail.com)
-- new behaviour: 8KB expandable to 64KB of internal RAM
--
-- MEMORY MAP
--    0000..1FFF : 8KB   8KB  block0 (upper 4KB used as DDR cache)
--    2000..3FFF : 8KB  16KB  block1 
--    4000..5FFF : 8KB  24KB  block2
--    6000..7FFF : 8KB  32KB  block3
--    8000..9FFF : 8KB  40KB  block4
--    A000..BFFF : 8KB  48KB  block5
--    C000..DFFF : 8KB  56KB  block6
--    E000..FFFF : 8KB  64KB  block7
---------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use work.mlite_pack.all;

library UNISIM;
use UNISIM.vcomponents.all;

entity boot_ram is
	generic(
		memory_type : string := "DEFAULT";
        --Number of 8KB blocks of internal RAM, up to 64KB (1 to 8)
        block_count : integer := 1
	); 
	port(
		clk               : in std_logic;
        enable            : in std_logic;
        write_byte_enable : in std_logic_vector(3 downto 0);
        address           : in std_logic_vector(31 downto 2);
        data_write        : in std_logic_vector(31 downto 0);
        data_read         : out std_logic_vector(31 downto 0)
	);
end; --entity boot_ram

architecture logic of boot_ram is
	--type
	type mem32_vector IS ARRAY (NATURAL RANGE<>) OF std_logic_vector(31 downto 0);

	--Which 8KB block
	alias block_sel: std_logic_vector(2 downto 0) is address(15 downto 13);

	--Address within a 8KB block (without lower two bits)
	alias block_addr : std_logic_vector(10 downto 0) is address(12 downto 2);

	--Block enable with 1 bit per memory block
	signal block_enable: std_logic_vector(7 downto 0);

	--Block Data Out
	signal block_do: mem32_vector(7 downto 0);

	--Remember which block was selected
	signal block_sel_buf: std_logic_vector(2 downto 0);

begin
	block_enable<= "00000001" when (enable='1') and (block_sel="000") else 
				   "00000010" when (enable='1') and (block_sel="001") else 
                   "00000100" when (enable='1') and (block_sel="010") else 
                   "00001000" when (enable='1') and (block_sel="011") else 
                   "00010000" when (enable='1') and (block_sel="100") else 
                   "00100000" when (enable='1') and (block_sel="101") else 
                   "01000000" when (enable='1') and (block_sel="110") else 
                   "10000000" when (enable='1') and (block_sel="111") else
                   "00000000";
  
	proc_blocksel: process (clk, block_sel) is
	begin
		if rising_edge(clk) then 
			block_sel_buf <= block_sel;
		end if;
	end process;

	proc_do: process (block_do, block_sel_buf) is
	begin
		data_read <= block_do(conv_integer(block_sel_buf));
	end process;
	
	-- BLOCKS generation
	block0: if (block_count > 0) generate
	begin

		ram_byte3 : RAMB16_S9
			generic map (
				INIT_00 => X"afafafafafafafafafafafafafafafaf2308000c241400ac273c243c243c273c",
				INIT_01 => X"8f8f8f8f8f8f8f8f8f8f8f8f8f8f8f8f8f230c008c8c3caf00af00af2340afaf",
				INIT_02 => X"acac0003373cac038cac8cac8cac8c243c000040034040033423038f038f8f8f",
				INIT_03 => X"00ac0300000034038c8c8c8c8c8c8c8c8c8c8c8c3403acacacacacacacacacac",
				INIT_04 => X"243c240caf3c00af2724033c2408a0100024241000283024a03c243c00000003",
				INIT_05 => X"afafaf3c2727038f8f02240c3c240c3c2408a01000242410002830022400a03c",
				INIT_06 => X"243c3c3c240c3c2412028c000200240002242400243c00240c3c1424a034afaf",
				INIT_07 => X"1200242410002832a2260c243c260c3c2408a0100024241000283202a2260c26",
				INIT_08 => X"afafafafafafaf272708248f8f8f8f8f3c00140008240c3c240c240c3c2608a2",
				INIT_09 => X"0c24240c240c0012001424142c2424142c2400142e24100010000c2424240000",
				INIT_0A => X"afafafafaf3caf2727038f8f8f8f8f8f028f240c240c00142a2602000c000826",
				INIT_0B => X"2727038f8f8f8f8f8f8fae16260c000800160014260c00a0028e3c3c003600af",
				INIT_0C => X"0c3c000c3c0c3c08000c3c0c00080014ae10000c020c24243c26afafafaf3caf",
				INIT_0D => X"31008cac001131008c001424083c24343c0003ac3c001030008c343c00000800",
				INIT_0E => X"001131008c2408001131008c00112c3000243c24343c00030014008024ac0011",
				INIT_0F => X"8c3c001030008c343c30038c343c0003ac3c241030008c343c00030014ac2424",
				INIT_10 => X"452e2e206b430a736461694a24038c3c0014ac00248c3c0824243c3c00000003",
				INIT_11 => X"000000000000000000006569612020740a004f3a63453a52006f202063746152",
				INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000"
			)
			port map (
				DO   => block_do(0)(31 downto 24), 
				DOP  => open, 
				ADDR => block_addr,
				CLK  => clk, 
				DI   => data_write(31 downto 24),
				DIP  => ZERO(0 downto 0),
				EN   => block_enable(0),
				SSR  => ZERO(0),
				WE   => write_byte_enable(3)
			);

		ram_byte2 : RAMB16_S9
			generic map (
				INIT_00 => X"b8afaeadacabaaa9a8a7a6a5a4a3a2a1bd000000a560a4a0bd1d8404a5059c1c",
				INIT_01 => X"b9b8afaeadacabaaa9a8a7a6a5a4a3a2a1a50086c6c406bb00bb00ba5a1abfb9",
				INIT_02 => X"919000405a1a06e0a606a606a606a6a505000084e0029b401bbd60bb60bbbabf",
				INIT_03 => X"00c4e0000085a2e09f9d9c9e979695949392919002e09f9d9c9e979695949392",
				INIT_04 => X"63038400bf0480b0bd42e00263006562c50606e004a7856340034202000000e0",
				INIT_05 => X"b2b3bf02bdbd20b0bf0084000484000442004446a40505e00387640042606002",
				INIT_06 => X"84100413840004423245d105470745444547520203040084000443424243b0b1",
				INIT_07 => X"1362030380124442203100840424001142004353830404a01165230060100073",
				INIT_08 => X"b2bfb0b1b3b4b5bdbd0084b0b1b2b3bf04024320008400040400840004100002",
				INIT_09 => X"0004040004002000405352606343526063434060435254205520001314150000",
				INIT_0A => X"bfb0b2b3b514b4bdbde0b0b1b2b3b4b520bf0400040020400210511100110010",
				INIT_0B => X"bdbde0b0b1b2b3b4b5bf4213100020002034204031000043b0431312009480b1",
				INIT_0C => X"0004200004000400200004002000205042512000600010111273bfb0b1b213b3",
				INIT_0D => X"0820a86620000820a8204706000307a50500e044022060632043420220200020",
				INIT_0E => X"20000820c8630020000820c82000686344070502c60620e02040208284622000",
				INIT_0F => X"42022060632043420242e042420220e043020360632043420220e04447a34263",
				INIT_10 => X"522e2e446968007364746e7542e042022044a0a34245030084420402202020e0",
				INIT_11 => X"020000401200400000000a6d7262666957004b207478206500726d4465206e3a",
				INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000"
			)
		port map (
			DO   => block_do(0)(23 downto 16),
			DOP  => open, 
			ADDR => block_addr,
			CLK  => clk, 
			DI   => data_write(23 downto 16),
			DIP  => ZERO(0 downto 0),
			EN   => block_enable(0),
			SSR  => ZERO(0),
			WE   => write_byte_enable(2)
		);
		
		ram_byte1 : RAMB16_S9
			generic map (
				INIT_00 => X"00000000000000000000000000000000ff00000100ff18000b000b0009008800",
				INIT_01 => X"000000000000000000000000000000000000012000002000d800d800ff700000",
				INIT_02 => X"0000000000100000000000000000000100000060006060000000000000000000",
				INIT_03 => X"0000002010000000000000000000000000000000000000000000000000000000",
				INIT_04 => X"0900080100008000ff090000ff00000028000000210000090000090000000000",
				INIT_05 => X"00000010ff00000000c8080100090100ff000000200000001900001809300000",
				INIT_06 => X"08000000080100000090002a903c00309000002e001010080100ff0000000000",
				INIT_07 => X"00100000009100000009010800090100ff000000180000008900001000090109",
				INIT_08 => X"00000000000000ff0001080000000000002eff08010801000001090100ff0000",
				INIT_09 => X"01000001000108009000ff0000ffff0000ff200000ff00080008010000008880",
				INIT_0A => X"00000000000000ff000000000000000010000001000108ff00008889018901ff",
				INIT_0B => X"ff00000000000000000009ff0001080108ff080000018800100900008086a800",
				INIT_0C => X"001008001001100108001001080108ff09000801200100000008000000000000",
				INIT_0D => X"0008000008ff00080008000001200000201000002008ff000800002008080108",
				INIT_0E => X"08ff000800000108ff0008000800000018ff20000020080008ff0800000008ff",
				INIT_0F => X"002008ff000800002000000000200800002000ff0008000020080018ff00ff00",
				INIT_10 => X"522e2e446e6500207220676d0000001008ff0028000010020908000008080800",
				INIT_11 => X"10000000101400000000006179696f6e61002100657000610079654473616e20",
				INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000"
			)
		port map (
			DO   => block_do(0)(15 downto 8),
			DOP  => open, 
			ADDR => block_addr,
			CLK  => clk, 
			DI   => data_write(15 downto 8),
			DIP  => ZERO(0 downto 0),
			EN   => block_enable(0),
			SSR  => ZERO(0),
			WE   => write_byte_enable(1)
		);

		ram_byte0 : RAMB16_S9
			generic map (
				INIT_00 => X"4c4844403c3834302c2824201c181410980e007f04fd2a00080020000000f001",
				INIT_01 => X"504c4844403c3834302c2824201c18141000e72410200060125c1058fc005450",
				INIT_02 => X"040000083c0048080c440840043c0068000000000800000801681360115c5854",
				INIT_03 => X"0c000810121900082c2824201c1814100c08040000082c2824201c1814100c08",
				INIT_04 => X"100050af14002110e8100800ff89000321303702020a0f170800100000000008",
				INIT_05 => X"1c202450d8180810142164af0010af00ffa5000321303702020a0f2117210800",
				INIT_06 => X"a00000007caf000435210000210002212101030078502168af00fd0100781418",
				INIT_07 => X"0321303702020a0f0810afa80010af00ffe5000321303702020a0f210817af10",
				INIT_08 => X"1c2c1418202428d028afb414181c20240000bf250b64af00fea410af00fff800",
				INIT_09 => X"a40820a408a42508210ca90e1a9fc9121abf21160ad020252225f7080d0a2121",
				INIT_0A => X"2c141c20280124d0300814181c202428212c0aa40da425dc10012100a40247ff",
				INIT_0B => X"d8300814181c2024282c00f101f7257625fb250501f221002100200021a02118",
				INIT_0C => X"970825bb0058009f25bb0058259a25f9000525f721afff3c00bc2414181c0020",
				INIT_0D => X"0225000025fc02250025070dc4000a20002108000025fc022500200025258a25",
				INIT_0E => X"25fc02250030e125fc02250025080a0f06fc001c2000250825ee2500010025fc",
				INIT_0F => X"000025fc012500200001080020002508000049fc0225002000250806ec00fc57",
				INIT_10 => X"4f002e5267630000656120708408000025fb00210400000e00e0000025252508",
				INIT_11 => X"001010200000207000000067206e726769000a006465006400216d5273636f43",
				INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000"
			)
		port map (
			DO   => block_do(0)(7 downto 0),
			DOP  => open, 
			ADDR => block_addr,
			CLK  => clk, 
			DI   => data_write(7 downto 0),
			DIP  => ZERO(0 downto 0),
			EN   => block_enable(0),
			SSR  => ZERO(0),
			WE   => write_byte_enable(0)
		);
		end generate; --block0
		

		block1: if (block_count > 1) generate
		begin

		ram_byte3 : RAMB16_S9
			generic map (
				INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000"
			)
			port map (
				DO   => block_do(1)(31 downto 24), 
				DOP  => open, 
				ADDR => block_addr,
				CLK  => clk, 
				DI   => data_write(31 downto 24),
				DIP  => ZERO(0 downto 0),
				EN   => block_enable(1),
				SSR  => ZERO(0),
				WE   => write_byte_enable(3)
			);

		ram_byte2 : RAMB16_S9
			generic map (
				INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000"
			)
			port map (
				DO   => block_do(1)(23 downto 16),
				DOP  => open, 
				ADDR => block_addr,
				CLK  => clk, 
				DI   => data_write(23 downto 16),
				DIP  => ZERO(0 downto 0),
				EN   => block_enable(1),
				SSR  => ZERO(0),
				WE   => write_byte_enable(2)
			);
		
		ram_byte1 : RAMB16_S9
			generic map (
			INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000"
		)
		port map (
		  DO   => block_do(1)(15 downto 8),
		  DOP  => open, 
		  ADDR => block_addr,
		  CLK  => clk, 
		  DI   => data_write(15 downto 8),
		  DIP  => ZERO(0 downto 0),
		  EN   => block_enable(1),
		  SSR  => ZERO(0),
		  WE   => write_byte_enable(1));

		ram_byte0 : RAMB16_S9
			generic map (
			INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000"
		)
		port map (
			DO   => block_do(1)(7 downto 0),
			DOP  => open, 
			ADDR => block_addr,
			CLK  => clk, 
			DI   => data_write(7 downto 0),
			DIP  => ZERO(0 downto 0),
			EN   => block_enable(1),
			SSR  => ZERO(0),
			WE   => write_byte_enable(0)
		);
		
	end generate; --block1
-- -------------------------------------------------------------------------------------------------------	
	block2: if (block_count > 2) generate
	begin

		ram_byte3 : RAMB16_S9
			generic map (
				INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000"
			)
			port map (
				DO   => block_do(2)(31 downto 24), 
				DOP  => open, 
				ADDR => block_addr,
				CLK  => clk, 
				DI   => data_write(31 downto 24),
				DIP  => ZERO(0 downto 0),
				EN   => block_enable(2),
				SSR  => ZERO(0),
				WE   => write_byte_enable(3)
			);

		ram_byte2 : RAMB16_S9
			generic map (
				INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000"
			)
			port map (
				DO   => block_do(2)(23 downto 16),
				DOP  => open, 
				ADDR => block_addr,
				CLK  => clk, 
				DI   => data_write(23 downto 16),
				DIP  => ZERO(0 downto 0),
				EN   => block_enable(2),
				SSR  => ZERO(0),
				WE   => write_byte_enable(2)
			);
	
		ram_byte1 : RAMB16_S9
			generic map (
				INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000"
			)
			port map (
				DO   => block_do(2)(15 downto 8),
				DOP  => open, 
				ADDR => block_addr,
				CLK  => clk, 
				DI   => data_write(15 downto 8),
				DIP  => ZERO(0 downto 0),
				EN   => block_enable(2),
				SSR  => ZERO(0),
				WE   => write_byte_enable(1)
			);

		ram_byte0 : RAMB16_S9
			generic map (
				INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000"
			)
		port map (
			DO   => block_do(2)(7 downto 0),
			DOP  => open, 
			ADDR => block_addr,
			CLK  => clk, 
			DI   => data_write(7 downto 0),
			DIP  => ZERO(0 downto 0),
			EN   => block_enable(2),
			SSR  => ZERO(0),
			WE   => write_byte_enable(0)
		);
		
	end generate; --block2
	
-- -------------------------------------------------------------------------------------------------------

	block3: if (block_count > 3) generate
	begin

		ram_byte3 : RAMB16_S9
			generic map (
				INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000"
			)
		port map (
			DO   => block_do(3)(31 downto 24), 
			DOP  => open, 
			ADDR => block_addr,
			CLK  => clk, 
			DI   => data_write(31 downto 24),
			DIP  => ZERO(0 downto 0),
			EN   => block_enable(3),
			SSR  => ZERO(0),
			WE   => write_byte_enable(3)
		);

    ram_byte2 : RAMB16_S9
		generic map (
			INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000"
		)
		port map (
			DO   => block_do(3)(23 downto 16),
			DOP  => open, 
			ADDR => block_addr,
			CLK  => clk, 
			DI   => data_write(23 downto 16),
			DIP  => ZERO(0 downto 0),
			EN   => block_enable(3),
			SSR  => ZERO(0),
			WE   => write_byte_enable(2)
		);
	
    ram_byte1 : RAMB16_S9
		generic map (
			INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000"
		)
		port map (
			DO   => block_do(3)(15 downto 8),
			DOP  => open, 
			ADDR => block_addr,
			CLK  => clk, 
			DI   => data_write(15 downto 8),
			DIP  => ZERO(0 downto 0),
			EN   => block_enable(3),
			SSR  => ZERO(0),
			WE   => write_byte_enable(1)
		);

    ram_byte0 : RAMB16_S9
		generic map (
			INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000"
		)
		port map (
			DO   => block_do(3)(7 downto 0),
			DOP  => open, 
			ADDR => block_addr,
			CLK  => clk, 
			DI   => data_write(7 downto 0),
			DIP  => ZERO(0 downto 0),
			EN   => block_enable(3),
			SSR  => ZERO(0),
			WE   => write_byte_enable(0)
		);
		
	end generate; --block3

-- -------------------------------------------------------------------------------------------------------

	block4: if (block_count > 4) generate
	begin

		ram_byte3 : RAMB16_S9
			generic map (
				INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000"
			)
			port map (
				DO   => block_do(4)(31 downto 24), 
				DOP  => open, 
				ADDR => block_addr,
				CLK  => clk, 
				DI   => data_write(31 downto 24),
				DIP  => ZERO(0 downto 0),
				EN   => block_enable(4),
				SSR  => ZERO(0),
				WE   => write_byte_enable(3)
			);

		ram_byte2 : RAMB16_S9
			generic map (
				INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000"
			)
			port map (
				DO   => block_do(4)(23 downto 16),
				DOP  => open, 
				ADDR => block_addr,
				CLK  => clk, 
				DI   => data_write(23 downto 16),
				DIP  => ZERO(0 downto 0),
				EN   => block_enable(4),
				SSR  => ZERO(0),
				WE   => write_byte_enable(2)
			);
	
		ram_byte1 : RAMB16_S9
			generic map (
				INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000"
			)
			port map (
				DO   => block_do(4)(15 downto 8),
				DOP  => open, 
				ADDR => block_addr,
				CLK  => clk, 
				DI   => data_write(15 downto 8),
				DIP  => ZERO(0 downto 0),
				EN   => block_enable(4),
				SSR  => ZERO(0),
				WE   => write_byte_enable(1)
			);

		ram_byte0 : RAMB16_S9
			generic map (
				INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000"
			)
			port map (
				DO   => block_do(4)(7 downto 0),
				DOP  => open, 
				ADDR => block_addr,
				CLK  => clk, 
				DI   => data_write(7 downto 0),
				DIP  => ZERO(0 downto 0),
				EN   => block_enable(4),
				SSR  => ZERO(0),
				WE   => write_byte_enable(0)
			);
		
   end generate; --block4

-- -------------------------------------------------------------------------------------------------------

	block5: if (block_count > 5) generate
	begin

    ram_byte3 : RAMB16_S9
   generic map (
INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000"
)
    port map (
      DO   => block_do(5)(31 downto 24), 
      DOP  => open, 
      ADDR => block_addr,
      CLK  => clk, 
      DI   => data_write(31 downto 24),
      DIP  => ZERO(0 downto 0),
      EN   => block_enable(5),
      SSR  => ZERO(0),
      WE   => write_byte_enable(3));

    ram_byte2 : RAMB16_S9
   generic map (
INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000"
)
    port map (
      DO   => block_do(5)(23 downto 16),
      DOP  => open, 
      ADDR => block_addr,
      CLK  => clk, 
      DI   => data_write(23 downto 16),
      DIP  => ZERO(0 downto 0),
      EN   => block_enable(5),
      SSR  => ZERO(0),
      WE   => write_byte_enable(2));
	
    ram_byte1 : RAMB16_S9
   generic map (
INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000"
)
    port map (
      DO   => block_do(5)(15 downto 8),
      DOP  => open, 
      ADDR => block_addr,
      CLK  => clk, 
      DI   => data_write(15 downto 8),
      DIP  => ZERO(0 downto 0),
      EN   => block_enable(5),
      SSR  => ZERO(0),
      WE   => write_byte_enable(1));

    ram_byte0 : RAMB16_S9
   generic map (
INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000"
)
    port map (
      DO   => block_do(5)(7 downto 0),
      DOP  => open, 
      ADDR => block_addr,
      CLK  => clk, 
      DI   => data_write(7 downto 0),
      DIP  => ZERO(0 downto 0),
      EN   => block_enable(5),
      SSR  => ZERO(0),
      WE   => write_byte_enable(0));
		
   end generate; --block5


   block6: if (block_count > 6) generate
	begin

    ram_byte3 : RAMB16_S9
   generic map (
INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000"
)
    port map (
      DO   => block_do(6)(31 downto 24), 
      DOP  => open, 
      ADDR => block_addr,
      CLK  => clk, 
      DI   => data_write(31 downto 24),
      DIP  => ZERO(0 downto 0),
      EN   => block_enable(6),
      SSR  => ZERO(0),
      WE   => write_byte_enable(3));

    ram_byte2 : RAMB16_S9
   generic map (
INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000"
)
    port map (
      DO   => block_do(6)(23 downto 16),
      DOP  => open, 
      ADDR => block_addr,
      CLK  => clk, 
      DI   => data_write(23 downto 16),
      DIP  => ZERO(0 downto 0),
      EN   => block_enable(6),
      SSR  => ZERO(0),
      WE   => write_byte_enable(2));
	
    ram_byte1 : RAMB16_S9
   generic map (
INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000"
)
    port map (
      DO   => block_do(6)(15 downto 8),
      DOP  => open, 
      ADDR => block_addr,
      CLK  => clk, 
      DI   => data_write(15 downto 8),
      DIP  => ZERO(0 downto 0),
      EN   => block_enable(6),
      SSR  => ZERO(0),
      WE   => write_byte_enable(1));

    ram_byte0 : RAMB16_S9
   generic map (
INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000"
)
    port map (
      DO   => block_do(6)(7 downto 0),
      DOP  => open, 
      ADDR => block_addr,
      CLK  => clk, 
      DI   => data_write(7 downto 0),
      DIP  => ZERO(0 downto 0),
      EN   => block_enable(6),
      SSR  => ZERO(0),
      WE   => write_byte_enable(0));
		
   end generate; --block6


   block7: if (block_count > 7) generate
	begin

    ram_byte3 : RAMB16_S9
   generic map (
INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000"
)
    port map (
      DO   => block_do(7)(31 downto 24), 
      DOP  => open, 
      ADDR => block_addr,
      CLK  => clk, 
      DI   => data_write(31 downto 24),
      DIP  => ZERO(0 downto 0),
      EN   => block_enable(7),
      SSR  => ZERO(0),
      WE   => write_byte_enable(3));

    ram_byte2 : RAMB16_S9
   generic map (
INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000"
)
    port map (
      DO   => block_do(7)(23 downto 16),
      DOP  => open, 
      ADDR => block_addr,
      CLK  => clk, 
      DI   => data_write(23 downto 16),
      DIP  => ZERO(0 downto 0),
      EN   => block_enable(7),
      SSR  => ZERO(0),
      WE   => write_byte_enable(2));
	
    ram_byte1 : RAMB16_S9
   generic map (
INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000"
)
    port map (
      DO   => block_do(7)(15 downto 8),
      DOP  => open, 
      ADDR => block_addr,
      CLK  => clk, 
      DI   => data_write(15 downto 8),
      DIP  => ZERO(0 downto 0),
      EN   => block_enable(7),
      SSR  => ZERO(0),
      WE   => write_byte_enable(1));

    ram_byte0 : RAMB16_S9
   generic map (
INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000"
)
    port map (
      DO   => block_do(7)(7 downto 0),
      DOP  => open, 
      ADDR => block_addr,
      CLK  => clk, 
      DI   => data_write(7 downto 0),
      DIP  => ZERO(0 downto 0),
      EN   => block_enable(7),
      SSR  => ZERO(0),
      WE   => write_byte_enable(0));
		
   end generate; --block7

end; --architecture logic
