library ieee;
use ieee.std_logic_1164.all;

entity dadda_mult is
	port(
		clk    : in  std_logic;
		rst    : in  std_logic;
		ce     : in  std_logic;
		sgn    : in  std_logic;
		a, b   : in  std_logic_vector(31 downto 0);
		c_mult : out std_logic_vector(63 downto 0)
	);
end;

architecture logic of dadda_mult is
	component full_adder
		port(
			a, b, c_in : in  std_logic;
			s, c_out   : out std_logic
		);
	end component;

	component half_adder
		port(
			a, b     : in  std_logic;
			s, c_out : out std_logic
		);
	end component;

	component flip_flop
		port(
			clk, rst : in  std_logic;
			ce, d    : in  std_logic;
			q        : out std_logic
		);
	end component;
	
	signal pp0, p0 : std_logic_vector(31 downto 0);
	signal pp1, p1 : std_logic_vector(31 downto 0);
	signal pp2, p2 : std_logic_vector(31 downto 0);
	signal pp3, p3 : std_logic_vector(31 downto 0);
	signal pp4, p4 : std_logic_vector(31 downto 0);
	signal pp5, p5 : std_logic_vector(31 downto 0);
	signal pp6, p6 : std_logic_vector(31 downto 0);
	signal pp7, p7 : std_logic_vector(31 downto 0);
	signal pp8, p8 : std_logic_vector(31 downto 0);
	signal pp9, p9 : std_logic_vector(31 downto 0);
	signal pp10, p10 : std_logic_vector(31 downto 0);
	signal pp11, p11 : std_logic_vector(31 downto 0);
	signal pp12, p12 : std_logic_vector(31 downto 0);
	signal pp13, p13 : std_logic_vector(31 downto 0);
	signal pp14, p14 : std_logic_vector(31 downto 0);
	signal pp15, p15 : std_logic_vector(31 downto 0);
	signal pp16, p16 : std_logic_vector(31 downto 0);
	signal pp17, p17 : std_logic_vector(31 downto 0);
	signal pp18, p18 : std_logic_vector(31 downto 0);
	signal pp19, p19 : std_logic_vector(31 downto 0);
	signal pp20, p20 : std_logic_vector(31 downto 0);
	signal pp21, p21 : std_logic_vector(31 downto 0);
	signal pp22, p22 : std_logic_vector(31 downto 0);
	signal pp23, p23 : std_logic_vector(31 downto 0);
	signal pp24, p24 : std_logic_vector(31 downto 0);
	signal pp25, p25 : std_logic_vector(31 downto 0);
	signal pp26, p26 : std_logic_vector(31 downto 0);
	signal pp27, p27 : std_logic_vector(31 downto 0);
	signal pp28, p28 : std_logic_vector(31 downto 0);
	signal pp29, p29 : std_logic_vector(31 downto 0);
	signal pp30, p30 : std_logic_vector(31 downto 0);
	signal pp31, p31 : std_logic_vector(31 downto 0);

	signal c297, s57, s56, s55, s54, s53, s52, s51, s50, s59, s58 : std_logic;
	signal c642, f119, c747, f114, f115, f116, f117, f110, f111, f112, f113 : std_logic;
	signal c745, c668, s196, c527, s159, c523, c899, c892, c893, c890, s850 : std_logic;
	signal c896, c897, c894, c895, c868, s583, c966, c967, c964, s829, s799 : std_logic;
	signal s798, c960, c961, s795, s794, s797, s796, s791, s790, s793, c864 : std_logic;
	signal c117, c444, c447, s249, s248, s243, s242, s241, s240, s247, s246 : std_logic;
	signal s245, s244, s965, c443, c442, f18, c709, s960, c702, c703, c700 : std_logic;
	signal c701, c706, c707, c704, c705, s308, s309, s306, s307, s304, s305 : std_logic;
	signal s303, s300, s301, c638, c639, c636, c637, c634, c635, c632, c633 : std_logic;
	signal c630, c631, c140, c141, c142, c143, c144, c145, c146, c147, c148 : std_logic;
	signal c149, c418, c419, c386, c387, c384, c385, c382, c383, c380, c381 : std_logic;
	signal c388, c590, c597, c562, c563, c561, c566, c567, c564, c568, c569 : std_logic;
	signal s461, f118, s878, s870, s871, s872, s874, s875, s876, s877, f40 : std_logic;
	signal f43, f42, f45, f44, f47, f46, f49, s625, s904, s905, s906 : std_logic;
	signal s907, s900, s901, s902, s903, s908, s909, s44, s45, s46, s47 : std_logic;
	signal s40, s41, s42, s43, s48, s49, c237, s379, f109, f108, f107 : std_logic;
	signal f106, f105, f104, c643, f102, f101, f100, c647, c39, c38, c646 : std_logic;
	signal c35, c34, c36, c31, c30, c33, c32, c644, s499, s496, s497 : std_logic;
	signal s494, s495, s492, s490, s491, c885, c884, c887, s658, c883, c882 : std_logic;
	signal c641, s655, s656, c640, s650, s651, s652, s653, s899, c971, c970 : std_logic;
	signal c973, c972, c975, c974, c977, c976, c979, c978, s180, s276, s277 : std_logic;
	signal s274, s217, s272, s273, s270, s278, s474, s475, s476, s477, s470 : std_logic;
	signal s471, s472, s473, s478, s479, s826, s318, s311, s310, s313, s315 : std_logic;
	signal s314, s317, s316, c629, c628, c621, c620, c623, c622, c625, c624 : std_logic;
	signal c627, c626, c153, c152, c151, c150, c157, c156, c155, c154, c409 : std_logic;
	signal s31, c159, c158, c898, c391, c390, c393, c392, c395, c394, c397 : std_logic;
	signal c396, c398, s828, c715, c714, c717, c711, c710, c713, c712, c719 : std_logic;
	signal c891, c579, c578, c575, c574, c577, c576, c570, c573, c572, c840 : std_logic;
	signal s869, s868, s863, s862, s861, s860, s867, s866, s865, s864, c843 : std_logic;
	signal s702, f56, f57, f54, f55, f52, f53, f51, f58, f59, s613 : std_logic;
	signal s917, s916, s915, s914, s913, s912, s910, c689, s919, s918, c654 : std_logic;
	signal s79, s78, c408, s71, s70, s73, s72, s75, s74, s77, s76 : std_logic;
	signal c656, s93, s92, s91, s90, s97, s96, s95, s94, s99, s98 : std_logic;
	signal c22, c23, c20, c26, c27, c24, c25, c28, c29, c657, s489 : std_logic;
	signal s481, s482, s485, s484, s487, s486, s649, s648, s647, s646, s645 : std_logic;
	signal s644, s643, s642, s641, s640, c488, s418, c765, c965, c962, c963 : std_logic;
	signal s873, c988, c989, c984, c985, c986, c987, c980, c981, c982, c983 : std_logic;
	signal c486, s261, s260, s263, s262, s265, s264, s267, s266, s269, s268 : std_logic;
	signal s792, s467, s466, s465, s464, s463, s462, s460, s469, s468, c804 : std_logic;
	signal c806, c802, c168, c169, c166, c167, c164, c165, c162, c163, c160 : std_logic;
	signal c161, c368, c369, c364, c365, c366, c367, c360, c361, c362, c363 : std_logic;
	signal c503, c760, c761, c762, c763, c764, c506, c766, c767, c768, c769 : std_logic;
	signal c508, c509, c500, c501, c502, c504, c505, c507, s108, s109, s104 : std_logic;
	signal s105, s106, s107, s100, s101, s102, s103, s610, c92, s612, c214 : std_logic;
	signal c215, c217, c210, c211, c212, c213, s936, s614, c218, s615, c184 : std_logic;
	signal c185, c186, c180, c181, c182, c183, s617, c189, s753, s922, s923 : std_logic;
	signal s920, c98, s927, s924, s925, s928, s929, s856, s857, s854, s852 : std_logic;
	signal s853, s68, s69, s66, s67, s65, s62, s63, s60, s61, f125 : std_logic;
	signal f124, s735, f120, f123, f122, s80, s81, s82, s83, s84, s85 : std_logic;
	signal s86, s87, s88, s89, c56, c55, c54, c53, c52, c51, c50 : std_logic;
	signal c59, c58, s678, s679, c851, s672, s673, s670, s671, s676, s677 : std_logic;
	signal s675, s805, c880, s631, s581, s582, s584, s585, s586, s587, s588 : std_logic;
	signal s589, c708, c991, c338, s298, s299, s294, s296, s297, s290, s291 : std_logic;
	signal s292, s293, s452, s453, s450, s451, s456, s454, s455, s458, s459 : std_logic;
	signal c188, s921, s302, s989, s926, c179, c178, c171, c170, c173, c172 : std_logic;
	signal c175, c174, c177, c176, c379, c378, c377, c376, c375, c374, c373 : std_logic;
	signal c372, c371, c370, c773, c772, c771, c770, c777, s199, c775, s198 : std_logic;
	signal c519, c513, c512, c511, c510, c517, c515, c514, s119, s118, s117 : std_logic;
	signal s116, s115, s114, s113, s112, s111, s110, s10, c819, c207, c205 : std_logic;
	signal c204, c203, c202, c200, c209, c208, c196, c195, c194, c193, c192 : std_logic;
	signal c191, c190, c199, c198, s681, c416, s939, s938, c417, s935, s934 : std_logic;
	signal s937, s931, c414, s933, s932, c415, c412, s684, c413, c410, c411 : std_logic;
	signal s841, s840, s843, s842, s845, s844, s847, s846, s849, c44, c45 : std_logic;
	signal c46, c47, c40, c41, c42, c43, c48, c49, s726, c799, c798 : std_logic;
	signal s665, s667, s666, c518, s660, s663, s662, s668, c795, s9, s8 : std_logic;
	signal s3, s1, s0, s7, s5, s4, s855, c389, s592, s591, s590 : std_logic;
	signal s597, s596, s595, c457, s599, s598, s721, f38, s394, s399, s858 : std_logic;
	signal s859, f90, s288, s287, s286, s285, s284, s283, s282, s281, s280 : std_logic;
	signal s449, s448, s445, s444, s447, s446, s441, s440, s443, s442, c834 : std_logic;
	signal c835, c836, c837, c830, c831, c833, s819, c839, f96, f97, c969 : std_logic;
	signal c953, c698, c699, c348, c349, c342, s6, c340, c341, c347, c344 : std_logic;
	signal c345, c824, c748, c749, c746, c744, c742, c743, c740, c741, c526 : std_logic;
	signal c57, c524, c525, c522, c520, c521, c528, c529, s128, s129, s122 : std_logic;
	signal s123, s120, s121, s126, s127, s124, s125, c828, c957, c232, c233 : std_logic;
	signal c230, c231, c236, c234, c238, c239, f89, f88, f85, f84, f87 : std_logic;
	signal f86, f81, f80, f83, f82, s948, s949, s940, s941, s942, s943 : std_logic;
	signal s944, s945, s946, s947, s773, c79, c78, c71, c70, c73, c72 : std_logic;
	signal c75, c74, c77, c76, c93, c91, c90, c97, c96, c95, c94 : std_logic;
	signal s618, s619, c99, s543, s822, s961, s879, s728, s729, s724, s725 : std_logic;
	signal s727, s720, s722, s723, s674, s438, s439, s430, s431, s432, s433 : std_logic;
	signal s434, s435, s436, s437, c827, c826, c825, c823, c822, c821, c820 : std_logic;
	signal c829, s544, s545, s546, s547, s540, s541, s542, s548, s549, c724 : std_logic;
	signal c355, c354, c357, c356, c351, c350, c353, c352, c359, c358, c688 : std_logic;
	signal c683, c682, c681, c680, c687, c686, c685, c759, f48, c751, c750 : std_logic;
	signal c753, c752, c755, c754, c757, c756, c530, c533, c532, c535, c537 : std_logic;
	signal c536, c539, c538, s135, s137, s136, s131, s130, s133, s132, s139 : std_logic;
	signal s138, s851, c684, f93, f91, c228, f94, f95, c225, c224, c227 : std_logic;
	signal c221, c220, c223, c222, s959, s958, s953, s952, s951, s950, s957 : std_logic;
	signal s956, s955, s954, f99, c758, c614, c947, c68, c69, c66, c67 : std_logic;
	signal c64, c65, c62, c63, c60, c61, c432, c80, c81, c82, c83 : std_logic;
	signal c84, c85, c86, c87, c89, s609, s608, c992, c433, c990, c534 : std_logic;
	signal c434, s830, c435, s739, s737, s736, s733, s732, s731, s730, c313 : std_logic;
	signal s134, c436, c430, c431, s833, s429, s428, s423, s422, s421, s420 : std_logic;
	signal s427, s426, s425, s424, c813, c810, c811, c816, c814, c437, s974 : std_logic;
	signal s557, s556, s555, s554, s553, s552, s551, s550, s559, s558, c320 : std_logic;
	signal c321, c322, c323, c324, c325, c326, c327, c328, c329, s295, c841 : std_logic;
	signal s140, s141, s142, s143, s144, s145, s146, s147, s148, s149, c788 : std_logic;
	signal c789, s386, s387, s384, s385, s382, s383, s381, s388, s389, c258 : std_logic;
	signal c250, c251, c252, c253, c254, c255, c256, c257, c922, f103, f9 : std_logic;
	signal f92, c546, s898, c547, s892, c229, s891, s896, s897, s894, s895 : std_logic;
	signal c678, c235, f98, c226, c548, c690, c445, c549, s966, s967, s964 : std_logic;
	signal s962, s963, c673, s968, s969, s638, s639, s636, s637, s634, s635 : std_logic;
	signal s632, s633, s630, c446, s714, c197, s708, s709, s703, s700, s701 : std_logic;
	signal s706, s707, s704, s705, c694, c441, c560, c695, c440, s493, s416 : std_logic;
	signal s417, s414, s415, s412, s413, s410, s411, s419, s201, c886, c809 : std_logic;
	signal c808, c805, c807, c691, c801, c800, c803, s659, s654, s209, s562 : std_logic;
	signal s563, s560, s561, s566, s567, s564, s565, c889, s568, s569, c888 : std_logic;
	signal c333, c332, c331, c330, c337, c336, c335, c334, c339, s508, f0 : std_logic;
	signal f1, f2, f3, f4, f5, f6, f7, f8, s153, s151, s150 : std_logic;
	signal s157, s156, s155, s154, c794, s158, c791, c790, c793, c792, s391 : std_logic;
	signal s390, s393, s392, s395, s397, s396, s398, c796, c206, c249, c248 : std_logic;
	signal c243, c242, c241, c240, c247, c246, c245, c244, c812, s885, s884 : std_logic;
	signal s887, s886, s881, s880, s883, c693, s888, c201, s971, s970, s973 : std_logic;
	signal s972, s975, s977, s976, s979, s978, s340, s628, s621, s620, s623 : std_logic;
	signal s622, s624, s627, s626, s344, s345, c817, c776, s715, s717, s716 : std_logic;
	signal s711, s710, s712, c774, s719, s718, c779, c782, c778, s401, s400 : std_logic;
	signal s403, s402, s405, s404, s407, s406, s409, s408, c780, c878, c879 : std_logic;
	signal c870, c871, c781, c873, c874, c875, c876, c877, c187, c293, c872 : std_logic;
	signal s579, s578, s575, s574, s576, s571, s570, s573, s572, c904, c905 : std_logic;
	signal c906, c900, c901, c902, c903, c456, c908, c909, c658, c659, c308 : std_logic;
	signal c309, c307, c304, c305, c302, c303, c300, c301, c458, c459, c516 : std_logic;
	signal c550, s168, s169, s166, s164, s165, s162, s163, s160, s161, s368 : std_logic;
	signal s369, s364, s365, s366, s360, s361, s362, s363, s275, c498, c499 : std_logic;
	signal c496, c497, c494, c495, c492, c493, c490, c491, c276, c277, c274 : std_logic;
	signal c275, c272, c273, c270, c271, s271, c278, c279, c475, c476, c477 : std_logic;
	signal c470, c471, c472, c473, s607, c478, c479, s606, s604, c584, s279 : std_logic;
	signal c216, c589, s184, s186, s187, s181, s182, s183, s188, s189, f23 : std_logic;
	signal f22, f21, c907, f27, f25, f24, s984, s985, f29, f28, s980 : std_logic;
	signal s982, s983, c37, s760, s761, s762, s763, s764, s766, s767, s768 : std_logic;
	signal s769, s577, f121, c306, c655, s890, c650, c651, c652, s483, c653 : std_logic;
	signal s319, c17, c869, c863, c862, c861, c860, c867, c866, c865, c219 : std_logic;
	signal s509, s312, s500, s501, s502, s503, s504, s505, s506, s507, c917 : std_logic;
	signal c916, c915, c914, c913, c912, c911, c910, c919, c918, c319, c318 : std_logic;
	signal c649, c648, c311, c310, c312, c315, c314, c317, c316, s214, s215 : std_logic;
	signal s216, s210, s211, s212, s213, s218, s219, s738, s179, s178, s171 : std_logic;
	signal s170, s173, s172, s175, s174, s177, s176, s734, s378, s377, s376 : std_logic;
	signal s375, s374, s373, s372, s371, s370, c489, c481, c480, c483, c482 : std_logic;
	signal c485, c484, c487, c261, c260, c263, c262, c265, c264, c267, c266 : std_logic;
	signal c269, c268, s930, c467, c466, c465, c464, c463, c462, c461, c460 : std_logic;
	signal c469, c468, c401, c474, c400, c718, c403, c402, c405, s629, c404 : std_logic;
	signal c407, c406, s752, s197, s195, s194, s193, s192, s191, s190, s19 : std_logic;
	signal s18, s13, s12, s11, s17, s16, s15, s14, c943, f30, f31 : std_logic;
	signal f32, f33, f34, f35, f36, f37, f39, s992, s991, s990, c399 : std_logic;
	signal s167, s772, s771, s770, s777, s776, s775, s774, s779, s778, s498 : std_logic;
	signal s848, s367, c856, c857, c854, c855, c852, c853, c850, c858, c859 : std_logic;
	signal c716, c21, f41, s519, s518, s513, s512, s511, s510, s517, s516 : std_logic;
	signal s515, s514, c923, c920, c921, c926, c927, c924, c925, c928, c929 : std_logic;
	signal c679, c672, c670, c671, c676, c677, c674, c675, s457, s207, s206 : std_logic;
	signal s205, s204, s203, s202, s200, s208, c815, c968, c818, s348, s349 : std_logic;
	signal s342, s343, s341, s346, s347, c298, c299, c294, c295, c296, c290 : std_logic;
	signal c291, c292, c452, c453, c450, c451, c108, c109, c454, c455, c104 : std_logic;
	signal c105, c106, c107, c100, c101, c102, c103, c571, c580, c581, c582 : std_logic;
	signal c583, c585, c586, c587, c588, c881, s834, s835, s836, s837, s831 : std_logic;
	signal s832, s664, c531, s838, s839, s657, s661, s746, s742, s669, s743 : std_logic;
	signal s740, s748, s749, s747, s744, s745, s741, s698, s699, c845, c844 : std_logic;
	signal c847, c846, s690, s691, s692, s693, s694, s695, s696, s697, s2 : std_logic;
	signal s526, s527, s524, s525, s522, s523, s520, s521, s528, s529, c939 : std_logic;
	signal c938, c935, c934, c937, c936, c931, c930, c933, c932, s580, s232 : std_logic;
	signal s233, s230, s231, s236, s234, s235, s238, s239, s593, s335, s355 : std_logic;
	signal s354, s357, s356, s351, s350, s353, s352, s359, s358, s185, s594 : std_logic;
	signal c665, c664, c667, c666, c661, c660, c663, c662, c669, c289, c288 : std_logic;
	signal c286, c285, c284, c283, c282, c281, c280, c449, c448, c119, c118 : std_logic;
	signal c116, c115, c114, c113, c112, c111, c110, c593, c592, c591, c596 : std_logic;
	signal c595, c594, c599, c598, s823, s911, c600, s827, s825, s824, s39 : std_logic;
	signal s38, s821, s820, s35, s34, s37, s36, s30, s33, s32, c842 : std_logic;
	signal c849, f19, s603, c848, f12, f13, f10, f11, f16, f17, f14 : std_logic;
	signal f15, s602, s601, s759, s758, s751, s750, s755, s754, s757, s756 : std_logic;
	signal s600, c783, c786, c787, c784, c785, s689, s688, s683, s682, s605 : std_logic;
	signal s680, s687, s686, s685, c426, f20, s988, f26, c343, s531, s530 : std_logic;
	signal s533, s532, s535, s534, s537, s536, s539, s538, s986, s987, s380 : std_logic;
	signal s981, c948, c949, c940, c941, c942, c944, c945, c946, s289, s229 : std_logic;
	signal s228, s225, s224, s227, s226, s221, s220, s223, s222, c728, c729 : std_logic;
	signal c725, c726, c727, c720, c721, c722, c723, s320, s321, s322, s323 : std_logic;
	signal s324, s325, s326, s327, s328, s329, c610, c611, c612, c613, c615 : std_logic;
	signal c616, c617, c618, c619, c438, c439, c128, c129, c122, c123, c120 : std_logic;
	signal c121, c126, c127, c124, c125, s765, c832, c287, c544, c545, c9 : std_logic;
	signal c8, c540, c541, c542, c543, c3, c2, c1, c0, c7, c6 : std_logic;
	signal c5, c4, c557, c88, c259, c838, s812, s813, s810, s811, s816 : std_logic;
	signal s817, s814, s815, s818, f69, f68, f67, f66, f65, f64, f63 : std_logic;
	signal f62, f61, f60, s22, s23, s20, s21, s26, s27, s24, s25 : std_logic;
	signal s28, s29, s611, s488, f50, c19, c18, s480, c13, c12, c11 : std_logic;
	signal c10, c16, c15, c14, s237, c645, s64, c565, s616, s782, s783 : std_logic;
	signal s780, s781, s786, s787, s784, s785, s788, s789, c959, c958, c952 : std_logic;
	signal c951, c950, c956, c955, c954, s801, s258, s259, s250, s251, s252 : std_logic;
	signal s253, s254, s255, s256, s257, c739, c738, c737, c736, c735, c734 : std_logic;
	signal c733, c732, c731, c730, s333, s332, s331, s330, s337, s336, s334 : std_logic;
	signal s339, s338, c797, s882, c603, c602, c601, c607, c606, c605, c604 : std_logic;
	signal c609, c608, c135, c134, c137, c136, c131, c130, c133, c132, c139 : std_logic;
	signal c138, c429, c428, c423, c422, c421, c420, c427, c425, c424, s152 : std_logic;
	signal c556, c555, c554, c553, c552, c551, c692, c559, c558, c346, c696 : std_logic;
	signal c697, s889, s809, s808, s804, s807, s806, s800, s803, s802, s713 : std_logic;
	signal s893, f78, f79, f74, f75, f76, f77, f70, f71, f72, f73 : std_logic;

begin
	pp0 <= (pp0'range => a(0)) and b;
	pp1 <= (pp1'range => a(1)) and b;
	pp2 <= (pp2'range => a(2)) and b;
	pp3 <= (pp3'range => a(3)) and b;
	pp4 <= (pp4'range => a(4)) and b;
	pp5 <= (pp5'range => a(5)) and b;
	pp6 <= (pp6'range => a(6)) and b;
	pp7 <= (pp7'range => a(7)) and b;
	pp8 <= (pp8'range => a(8)) and b;
	pp9 <= (pp9'range => a(9)) and b;
	pp10 <= (pp10'range => a(10)) and b;
	pp11 <= (pp11'range => a(11)) and b;
	pp12 <= (pp12'range => a(12)) and b;
	pp13 <= (pp13'range => a(13)) and b;
	pp14 <= (pp14'range => a(14)) and b;
	pp15 <= (pp15'range => a(15)) and b;
	pp16 <= (pp16'range => a(16)) and b;
	pp17 <= (pp17'range => a(17)) and b;
	pp18 <= (pp18'range => a(18)) and b;
	pp19 <= (pp19'range => a(19)) and b;
	pp20 <= (pp20'range => a(20)) and b;
	pp21 <= (pp21'range => a(21)) and b;
	pp22 <= (pp22'range => a(22)) and b;
	pp23 <= (pp23'range => a(23)) and b;
	pp24 <= (pp24'range => a(24)) and b;
	pp25 <= (pp25'range => a(25)) and b;
	pp26 <= (pp26'range => a(26)) and b;
	pp27 <= (pp27'range => a(27)) and b;
	pp28 <= (pp28'range => a(28)) and b;
	pp29 <= (pp29'range => a(29)) and b;
	pp30 <= (pp30'range => a(30)) and b;
	pp31 <= (pp31'range => a(31)) and b;

	p0 <= pp0 when sgn = '0' else (not pp0(31)) & pp0(30 downto 0);
	p1 <= pp1 when sgn = '0' else (not pp1(31)) & pp1(30 downto 0);
	p2 <= pp2 when sgn = '0' else (not pp2(31)) & pp2(30 downto 0);
	p3 <= pp3 when sgn = '0' else (not pp3(31)) & pp3(30 downto 0);
	p4 <= pp4 when sgn = '0' else (not pp4(31)) & pp4(30 downto 0);
	p5 <= pp5 when sgn = '0' else (not pp5(31)) & pp5(30 downto 0);
	p6 <= pp6 when sgn = '0' else (not pp6(31)) & pp6(30 downto 0);
	p7 <= pp7 when sgn = '0' else (not pp7(31)) & pp7(30 downto 0);
	p8 <= pp8 when sgn = '0' else (not pp8(31)) & pp8(30 downto 0);
	p9 <= pp9 when sgn = '0' else (not pp9(31)) & pp9(30 downto 0);
	p10 <= pp10 when sgn = '0' else (not pp10(31)) & pp10(30 downto 0);
	p11 <= pp11 when sgn = '0' else (not pp11(31)) & pp11(30 downto 0);
	p12 <= pp12 when sgn = '0' else (not pp12(31)) & pp12(30 downto 0);
	p13 <= pp13 when sgn = '0' else (not pp13(31)) & pp13(30 downto 0);
	p14 <= pp14 when sgn = '0' else (not pp14(31)) & pp14(30 downto 0);
	p15 <= pp15 when sgn = '0' else (not pp15(31)) & pp15(30 downto 0);
	p16 <= pp16 when sgn = '0' else (not pp16(31)) & pp16(30 downto 0);
	p17 <= pp17 when sgn = '0' else (not pp17(31)) & pp17(30 downto 0);
	p18 <= pp18 when sgn = '0' else (not pp18(31)) & pp18(30 downto 0);
	p19 <= pp19 when sgn = '0' else (not pp19(31)) & pp19(30 downto 0);
	p20 <= pp20 when sgn = '0' else (not pp20(31)) & pp20(30 downto 0);
	p21 <= pp21 when sgn = '0' else (not pp21(31)) & pp21(30 downto 0);
	p22 <= pp22 when sgn = '0' else (not pp22(31)) & pp22(30 downto 0);
	p23 <= pp23 when sgn = '0' else (not pp23(31)) & pp23(30 downto 0);
	p24 <= pp24 when sgn = '0' else (not pp24(31)) & pp24(30 downto 0);
	p25 <= pp25 when sgn = '0' else (not pp25(31)) & pp25(30 downto 0);
	p26 <= pp26 when sgn = '0' else (not pp26(31)) & pp26(30 downto 0);
	p27 <= pp27 when sgn = '0' else (not pp27(31)) & pp27(30 downto 0);
	p28 <= pp28 when sgn = '0' else (not pp28(31)) & pp28(30 downto 0);
	p29 <= pp29 when sgn = '0' else (not pp29(31)) & pp29(30 downto 0);
	p30 <= pp30 when sgn = '0' else (not pp30(31)) & pp30(30 downto 0);
	p31 <= pp31 when sgn = '0' else pp31(31) & (not pp31(30 downto 0));

	adder0000: half_adder port map(a => p0(28), b => p1(27), s => s0, c_out => c0);
	adder0001: full_adder port map(a => p0(29), b => p1(28), c_in => c0, s => s1, c_out => c1);
	adder0002: half_adder port map(a => p2(27), b => p3(26), s => s2, c_out => c2);
	adder0003: full_adder port map(a => c1, b => p0(30), c_in => c2, s => s3, c_out => c3);
	adder0004: full_adder port map(a => p2(28), b => p3(27), c_in => p1(29), s => s4, c_out => c4);
	adder0005: half_adder port map(a => p4(26), b => p5(25), s => s5, c_out => c5);
	adder0006: full_adder port map(a => c4, b => c3, c_in => c5, s => s6, c_out => c6);
	adder0007: full_adder port map(a => p1(30), b => p2(29), c_in => p0(31), s => s7, c_out => c7);
	adder0008: full_adder port map(a => p4(27), b => p5(26), c_in => p3(28), s => s8, c_out => c8);
	adder0009: half_adder port map(a => p6(25), b => p7(24), s => s9, c_out => c9);
	adder0010: full_adder port map(a => c8, b => c7, c_in => c9, s => s10, c_out => c10);
	adder0011: full_adder port map(a => sgn, b => p1(31), c_in => c6, s => s11, c_out => c11);
	adder0012: full_adder port map(a => p3(29), b => p4(28), c_in => p2(30), s => s12, c_out => c12);
	adder0013: full_adder port map(a => p6(26), b => p7(25), c_in => p5(27), s => s13, c_out => c13);
	adder0014: full_adder port map(a => c12, b => c11, c_in => c13, s => s14, c_out => c14);
	adder0015: full_adder port map(a => p2(31), b => p3(30), c_in => c10, s => s15, c_out => c15);
	adder0016: full_adder port map(a => p5(28), b => p6(27), c_in => p4(29), s => s16, c_out => c16);
	adder0017: full_adder port map(a => c15, b => c14, c_in => c16, s => s17, c_out => c17);
	adder0018: full_adder port map(a => p4(30), b => p5(29), c_in => p3(31), s => s18, c_out => c18);
	adder0019: full_adder port map(a => c17, b => p4(31), c_in => c18, s => s19, c_out => c19);
	adder0020: half_adder port map(a => p0(19), b => p1(18), s => s20, c_out => c20);
	adder0021: full_adder port map(a => p0(20), b => p1(19), c_in => c20, s => s21, c_out => c21);
	adder0022: half_adder port map(a => p2(18), b => p3(17), s => s22, c_out => c22);
	adder0023: full_adder port map(a => c21, b => p0(21), c_in => c22, s => s23, c_out => c23);
	adder0024: full_adder port map(a => p2(19), b => p3(18), c_in => p1(20), s => s24, c_out => c24);
	adder0025: half_adder port map(a => p4(17), b => p5(16), s => s25, c_out => c25);
	adder0026: full_adder port map(a => c24, b => c23, c_in => c25, s => s26, c_out => c26);
	adder0027: full_adder port map(a => p1(21), b => p2(20), c_in => p0(22), s => s27, c_out => c27);
	adder0028: full_adder port map(a => p4(18), b => p5(17), c_in => p3(19), s => s28, c_out => c28);
	adder0029: half_adder port map(a => p6(16), b => p7(15), s => s29, c_out => c29);
	adder0030: full_adder port map(a => c28, b => c27, c_in => c29, s => s30, c_out => c30);
	adder0031: full_adder port map(a => p0(23), b => p1(22), c_in => c26, s => s31, c_out => c31);
	adder0032: full_adder port map(a => p3(20), b => p4(19), c_in => p2(21), s => s32, c_out => c32);
	adder0033: full_adder port map(a => p6(17), b => p7(16), c_in => p5(18), s => s33, c_out => c33);
	adder0034: half_adder port map(a => p8(15), b => p9(14), s => s34, c_out => c34);
	adder0035: full_adder port map(a => c33, b => c32, c_in => c34, s => s35, c_out => c35);
	adder0036: full_adder port map(a => c30, b => p0(24), c_in => c31, s => s36, c_out => c36);
	adder0037: full_adder port map(a => p2(22), b => p3(21), c_in => p1(23), s => s37, c_out => c37);
	adder0038: full_adder port map(a => p5(19), b => p6(18), c_in => p4(20), s => s38, c_out => c38);
	adder0039: full_adder port map(a => p8(16), b => p9(15), c_in => p7(17), s => s39, c_out => c39);
	adder0040: half_adder port map(a => p10(14), b => p11(13), s => s40, c_out => c40);
	adder0041: full_adder port map(a => c39, b => c38, c_in => c40, s => s41, c_out => c41);
	adder0042: full_adder port map(a => c36, b => c35, c_in => c37, s => s42, c_out => c42);
	adder0043: full_adder port map(a => p1(24), b => p2(23), c_in => p0(25), s => s43, c_out => c43);
	adder0044: full_adder port map(a => p4(21), b => p5(20), c_in => p3(22), s => s44, c_out => c44);
	adder0045: full_adder port map(a => p7(18), b => p8(17), c_in => p6(19), s => s45, c_out => c45);
	adder0046: full_adder port map(a => p10(15), b => p11(14), c_in => p9(16), s => s46, c_out => c46);
	adder0047: half_adder port map(a => p12(13), b => p13(12), s => s47, c_out => c47);
	adder0048: full_adder port map(a => c46, b => c45, c_in => c47, s => s48, c_out => c48);
	adder0049: full_adder port map(a => c43, b => c42, c_in => c44, s => s49, c_out => c49);
	adder0050: full_adder port map(a => p0(26), b => p1(25), c_in => c41, s => s50, c_out => c50);
	adder0051: full_adder port map(a => p3(23), b => p4(22), c_in => p2(24), s => s51, c_out => c51);
	adder0052: full_adder port map(a => p6(20), b => p7(19), c_in => p5(21), s => s52, c_out => c52);
	adder0053: full_adder port map(a => p9(17), b => p10(16), c_in => p8(18), s => s53, c_out => c53);
	adder0054: full_adder port map(a => p12(14), b => p13(13), c_in => p11(15), s => s54, c_out => c54);
	adder0055: half_adder port map(a => p14(12), b => p15(11), s => s55, c_out => c55);
	adder0056: full_adder port map(a => c54, b => c53, c_in => c55, s => s56, c_out => c56);
	adder0057: full_adder port map(a => c51, b => c50, c_in => c52, s => s57, c_out => c57);
	adder0058: full_adder port map(a => c48, b => p0(27), c_in => c49, s => s58, c_out => c58);
	adder0059: full_adder port map(a => p2(25), b => p3(24), c_in => p1(26), s => s59, c_out => c59);
	adder0060: full_adder port map(a => p5(22), b => p6(21), c_in => p4(23), s => s60, c_out => c60);
	adder0061: full_adder port map(a => p8(19), b => p9(18), c_in => p7(20), s => s61, c_out => c61);
	adder0062: full_adder port map(a => p11(16), b => p12(15), c_in => p10(17), s => s62, c_out => c62);
	adder0063: full_adder port map(a => p14(13), b => p15(12), c_in => p13(14), s => s63, c_out => c63);
	adder0064: half_adder port map(a => p16(11), b => p17(10), s => s64, c_out => c64);
	adder0065: full_adder port map(a => c63, b => c62, c_in => c64, s => s65, c_out => c65);
	adder0066: full_adder port map(a => c60, b => c59, c_in => c61, s => s66, c_out => c66);
	adder0067: full_adder port map(a => c57, b => c56, c_in => c58, s => s67, c_out => c67);
	adder0068: full_adder port map(a => p3(25), b => p4(24), c_in => p2(26), s => s68, c_out => c68);
	adder0069: full_adder port map(a => p6(22), b => p7(21), c_in => p5(23), s => s69, c_out => c69);
	adder0070: full_adder port map(a => p9(19), b => p10(18), c_in => p8(20), s => s70, c_out => c70);
	adder0071: full_adder port map(a => p12(16), b => p13(15), c_in => p11(17), s => s71, c_out => c71);
	adder0072: full_adder port map(a => p15(13), b => p16(12), c_in => p14(14), s => s72, c_out => c72);
	adder0073: full_adder port map(a => p18(10), b => p19(9), c_in => p17(11), s => s73, c_out => c73);
	adder0074: full_adder port map(a => c72, b => c71, c_in => c73, s => s74, c_out => c74);
	adder0075: full_adder port map(a => c69, b => c68, c_in => c70, s => s75, c_out => c75);
	adder0076: full_adder port map(a => c66, b => c65, c_in => c67, s => s76, c_out => c76);
	adder0077: full_adder port map(a => p5(24), b => p6(23), c_in => p4(25), s => s77, c_out => c77);
	adder0078: full_adder port map(a => p8(21), b => p9(20), c_in => p7(22), s => s78, c_out => c78);
	adder0079: full_adder port map(a => p11(18), b => p12(17), c_in => p10(19), s => s79, c_out => c79);
	adder0080: full_adder port map(a => p14(15), b => p15(14), c_in => p13(16), s => s80, c_out => c80);
	adder0081: full_adder port map(a => p17(12), b => p18(11), c_in => p16(13), s => s81, c_out => c81);
	adder0082: full_adder port map(a => p20(9), b => p21(8), c_in => p19(10), s => s82, c_out => c82);
	adder0083: full_adder port map(a => c81, b => c80, c_in => c82, s => s83, c_out => c83);
	adder0084: full_adder port map(a => c78, b => c77, c_in => c79, s => s84, c_out => c84);
	adder0085: full_adder port map(a => c75, b => c74, c_in => c76, s => s85, c_out => c85);
	adder0086: full_adder port map(a => p7(23), b => p8(22), c_in => p6(24), s => s86, c_out => c86);
	adder0087: full_adder port map(a => p10(20), b => p11(19), c_in => p9(21), s => s87, c_out => c87);
	adder0088: full_adder port map(a => p13(17), b => p14(16), c_in => p12(18), s => s88, c_out => c88);
	adder0089: full_adder port map(a => p16(14), b => p17(13), c_in => p15(15), s => s89, c_out => c89);
	adder0090: full_adder port map(a => p19(11), b => p20(10), c_in => p18(12), s => s90, c_out => c90);
	adder0091: full_adder port map(a => p22(8), b => p23(7), c_in => p21(9), s => s91, c_out => c91);
	adder0092: full_adder port map(a => c90, b => c89, c_in => c91, s => s92, c_out => c92);
	adder0093: full_adder port map(a => c87, b => c86, c_in => c88, s => s93, c_out => c93);
	adder0094: full_adder port map(a => c84, b => c83, c_in => c85, s => s94, c_out => c94);
	adder0095: full_adder port map(a => p9(22), b => p10(21), c_in => p8(23), s => s95, c_out => c95);
	adder0096: full_adder port map(a => p12(19), b => p13(18), c_in => p11(20), s => s96, c_out => c96);
	adder0097: full_adder port map(a => p15(16), b => p16(15), c_in => p14(17), s => s97, c_out => c97);
	adder0098: full_adder port map(a => p18(13), b => p19(12), c_in => p17(14), s => s98, c_out => c98);
	adder0099: full_adder port map(a => p21(10), b => p22(9), c_in => p20(11), s => s99, c_out => c99);
	adder0100: full_adder port map(a => p24(7), b => p25(6), c_in => p23(8), s => s100, c_out => c100);
	adder0101: full_adder port map(a => c99, b => c98, c_in => c100, s => s101, c_out => c101);
	adder0102: full_adder port map(a => c96, b => c95, c_in => c97, s => s102, c_out => c102);
	adder0103: full_adder port map(a => c93, b => c92, c_in => c94, s => s103, c_out => c103);
	adder0104: full_adder port map(a => p9(23), b => p10(22), c_in => p8(24), s => s104, c_out => c104);
	adder0105: full_adder port map(a => p12(20), b => p13(19), c_in => p11(21), s => s105, c_out => c105);
	adder0106: full_adder port map(a => p15(17), b => p16(16), c_in => p14(18), s => s106, c_out => c106);
	adder0107: full_adder port map(a => p18(14), b => p19(13), c_in => p17(15), s => s107, c_out => c107);
	adder0108: full_adder port map(a => p21(11), b => p22(10), c_in => p20(12), s => s108, c_out => c108);
	adder0109: full_adder port map(a => p24(8), b => p25(7), c_in => p23(9), s => s109, c_out => c109);
	adder0110: full_adder port map(a => c108, b => c107, c_in => c109, s => s110, c_out => c110);
	adder0111: full_adder port map(a => c105, b => c104, c_in => c106, s => s111, c_out => c111);
	adder0112: full_adder port map(a => c102, b => c101, c_in => c103, s => s112, c_out => c112);
	adder0113: full_adder port map(a => p8(25), b => p9(24), c_in => p7(26), s => s113, c_out => c113);
	adder0114: full_adder port map(a => p11(22), b => p12(21), c_in => p10(23), s => s114, c_out => c114);
	adder0115: full_adder port map(a => p14(19), b => p15(18), c_in => p13(20), s => s115, c_out => c115);
	adder0116: full_adder port map(a => p17(16), b => p18(15), c_in => p16(17), s => s116, c_out => c116);
	adder0117: full_adder port map(a => p20(13), b => p21(12), c_in => p19(14), s => s117, c_out => c117);
	adder0118: full_adder port map(a => p23(10), b => p24(9), c_in => p22(11), s => s118, c_out => c118);
	adder0119: full_adder port map(a => c117, b => c116, c_in => c118, s => s119, c_out => c119);
	adder0120: full_adder port map(a => c114, b => c113, c_in => c115, s => s120, c_out => c120);
	adder0121: full_adder port map(a => c111, b => c110, c_in => c112, s => s121, c_out => c121);
	adder0122: full_adder port map(a => p7(27), b => p8(26), c_in => p6(28), s => s122, c_out => c122);
	adder0123: full_adder port map(a => p10(24), b => p11(23), c_in => p9(25), s => s123, c_out => c123);
	adder0124: full_adder port map(a => p13(21), b => p14(20), c_in => p12(22), s => s124, c_out => c124);
	adder0125: full_adder port map(a => p16(18), b => p17(17), c_in => p15(19), s => s125, c_out => c125);
	adder0126: full_adder port map(a => p19(15), b => p20(14), c_in => p18(16), s => s126, c_out => c126);
	adder0127: full_adder port map(a => p22(12), b => p23(11), c_in => p21(13), s => s127, c_out => c127);
	adder0128: full_adder port map(a => c126, b => c125, c_in => c127, s => s128, c_out => c128);
	adder0129: full_adder port map(a => c123, b => c122, c_in => c124, s => s129, c_out => c129);
	adder0130: full_adder port map(a => c120, b => c119, c_in => c121, s => s130, c_out => c130);
	adder0131: full_adder port map(a => p6(29), b => p7(28), c_in => p5(30), s => s131, c_out => c131);
	adder0132: full_adder port map(a => p9(26), b => p10(25), c_in => p8(27), s => s132, c_out => c132);
	adder0133: full_adder port map(a => p12(23), b => p13(22), c_in => p11(24), s => s133, c_out => c133);
	adder0134: full_adder port map(a => p15(20), b => p16(19), c_in => p14(21), s => s134, c_out => c134);
	adder0135: full_adder port map(a => p18(17), b => p19(16), c_in => p17(18), s => s135, c_out => c135);
	adder0136: full_adder port map(a => p21(14), b => p22(13), c_in => p20(15), s => s136, c_out => c136);
	adder0137: full_adder port map(a => c135, b => c134, c_in => c136, s => s137, c_out => c137);
	adder0138: full_adder port map(a => c132, b => c131, c_in => c133, s => s138, c_out => c138);
	adder0139: full_adder port map(a => c129, b => c128, c_in => c130, s => s139, c_out => c139);
	adder0140: full_adder port map(a => p5(31), b => p6(30), c_in => c19, s => s140, c_out => c140);
	adder0141: full_adder port map(a => p8(28), b => p9(27), c_in => p7(29), s => s141, c_out => c141);
	adder0142: full_adder port map(a => p11(25), b => p12(24), c_in => p10(26), s => s142, c_out => c142);
	adder0143: full_adder port map(a => p14(22), b => p15(21), c_in => p13(23), s => s143, c_out => c143);
	adder0144: full_adder port map(a => p17(19), b => p18(18), c_in => p16(20), s => s144, c_out => c144);
	adder0145: full_adder port map(a => p20(16), b => p21(15), c_in => p19(17), s => s145, c_out => c145);
	adder0146: full_adder port map(a => c144, b => c143, c_in => c145, s => s146, c_out => c146);
	adder0147: full_adder port map(a => c141, b => c140, c_in => c142, s => s147, c_out => c147);
	adder0148: full_adder port map(a => c138, b => c137, c_in => c139, s => s148, c_out => c148);
	adder0149: full_adder port map(a => p7(30), b => p8(29), c_in => p6(31), s => s149, c_out => c149);
	adder0150: full_adder port map(a => p10(27), b => p11(26), c_in => p9(28), s => s150, c_out => c150);
	adder0151: full_adder port map(a => p13(24), b => p14(23), c_in => p12(25), s => s151, c_out => c151);
	adder0152: full_adder port map(a => p16(21), b => p17(20), c_in => p15(22), s => s152, c_out => c152);
	adder0153: full_adder port map(a => p19(18), b => p20(17), c_in => p18(19), s => s153, c_out => c153);
	adder0154: full_adder port map(a => c152, b => c151, c_in => c153, s => s154, c_out => c154);
	adder0155: full_adder port map(a => c149, b => c148, c_in => c150, s => s155, c_out => c155);
	adder0156: full_adder port map(a => c146, b => p7(31), c_in => c147, s => s156, c_out => c156);
	adder0157: full_adder port map(a => p9(29), b => p10(28), c_in => p8(30), s => s157, c_out => c157);
	adder0158: full_adder port map(a => p12(26), b => p13(25), c_in => p11(27), s => s158, c_out => c158);
	adder0159: full_adder port map(a => p15(23), b => p16(22), c_in => p14(24), s => s159, c_out => c159);
	adder0160: full_adder port map(a => p18(20), b => p19(19), c_in => p17(21), s => s160, c_out => c160);
	adder0161: full_adder port map(a => c159, b => c158, c_in => c160, s => s161, c_out => c161);
	adder0162: full_adder port map(a => c156, b => c155, c_in => c157, s => s162, c_out => c162);
	adder0163: full_adder port map(a => p8(31), b => p9(30), c_in => c154, s => s163, c_out => c163);
	adder0164: full_adder port map(a => p11(28), b => p12(27), c_in => p10(29), s => s164, c_out => c164);
	adder0165: full_adder port map(a => p14(25), b => p15(24), c_in => p13(26), s => s165, c_out => c165);
	adder0166: full_adder port map(a => p17(22), b => p18(21), c_in => p16(23), s => s166, c_out => c166);
	adder0167: full_adder port map(a => c165, b => c164, c_in => c166, s => s167, c_out => c167);
	adder0168: full_adder port map(a => c162, b => c161, c_in => c163, s => s168, c_out => c168);
	adder0169: full_adder port map(a => p10(30), b => p11(29), c_in => p9(31), s => s169, c_out => c169);
	adder0170: full_adder port map(a => p13(27), b => p14(26), c_in => p12(28), s => s170, c_out => c170);
	adder0171: full_adder port map(a => p16(24), b => p17(23), c_in => p15(25), s => s171, c_out => c171);
	adder0172: full_adder port map(a => c170, b => c169, c_in => c171, s => s172, c_out => c172);
	adder0173: full_adder port map(a => c167, b => p10(31), c_in => c168, s => s173, c_out => c173);
	adder0174: full_adder port map(a => p12(29), b => p13(28), c_in => p11(30), s => s174, c_out => c174);
	adder0175: full_adder port map(a => p15(26), b => p16(25), c_in => p14(27), s => s175, c_out => c175);
	adder0176: full_adder port map(a => c174, b => c173, c_in => c175, s => s176, c_out => c176);
	adder0177: full_adder port map(a => p11(31), b => p12(30), c_in => c172, s => s177, c_out => c177);
	adder0178: full_adder port map(a => p14(28), b => p15(27), c_in => p13(29), s => s178, c_out => c178);
	adder0179: full_adder port map(a => c177, b => c176, c_in => c178, s => s179, c_out => c179);
	adder0180: full_adder port map(a => p13(30), b => p14(29), c_in => p12(31), s => s180, c_out => c180);
	adder0181: full_adder port map(a => c179, b => p13(31), c_in => c180, s => s181, c_out => c181);
	adder0182: half_adder port map(a => p0(13), b => p1(12), s => s182, c_out => c182);
	adder0183: full_adder port map(a => p0(14), b => p1(13), c_in => c182, s => s183, c_out => c183);
	adder0184: half_adder port map(a => p2(12), b => p3(11), s => s184, c_out => c184);
	adder0185: full_adder port map(a => c183, b => p0(15), c_in => c184, s => s185, c_out => c185);
	adder0186: full_adder port map(a => p2(13), b => p3(12), c_in => p1(14), s => s186, c_out => c186);
	adder0187: half_adder port map(a => p4(11), b => p5(10), s => s187, c_out => c187);
	adder0188: full_adder port map(a => c186, b => c185, c_in => c187, s => s188, c_out => c188);
	adder0189: full_adder port map(a => p1(15), b => p2(14), c_in => p0(16), s => s189, c_out => c189);
	adder0190: full_adder port map(a => p4(12), b => p5(11), c_in => p3(13), s => s190, c_out => c190);
	adder0191: half_adder port map(a => p6(10), b => p7(9), s => s191, c_out => c191);
	adder0192: full_adder port map(a => c190, b => c189, c_in => c191, s => s192, c_out => c192);
	adder0193: full_adder port map(a => p0(17), b => p1(16), c_in => c188, s => s193, c_out => c193);
	adder0194: full_adder port map(a => p3(14), b => p4(13), c_in => p2(15), s => s194, c_out => c194);
	adder0195: full_adder port map(a => p6(11), b => p7(10), c_in => p5(12), s => s195, c_out => c195);
	adder0196: half_adder port map(a => p8(9), b => p9(8), s => s196, c_out => c196);
	adder0197: full_adder port map(a => c195, b => c194, c_in => c196, s => s197, c_out => c197);
	adder0198: full_adder port map(a => c192, b => p0(18), c_in => c193, s => s198, c_out => c198);
	adder0199: full_adder port map(a => p2(16), b => p3(15), c_in => p1(17), s => s199, c_out => c199);
	adder0200: full_adder port map(a => p5(13), b => p6(12), c_in => p4(14), s => s200, c_out => c200);
	adder0201: full_adder port map(a => p8(10), b => p9(9), c_in => p7(11), s => s201, c_out => c201);
	adder0202: half_adder port map(a => p10(8), b => p11(7), s => s202, c_out => c202);
	adder0203: full_adder port map(a => c201, b => c200, c_in => c202, s => s203, c_out => c203);
	adder0204: full_adder port map(a => c198, b => c197, c_in => c199, s => s204, c_out => c204);
	adder0205: full_adder port map(a => p3(16), b => p4(15), c_in => p2(17), s => s205, c_out => c205);
	adder0206: full_adder port map(a => p6(13), b => p7(12), c_in => p5(14), s => s206, c_out => c206);
	adder0207: full_adder port map(a => p9(10), b => p10(9), c_in => p8(11), s => s207, c_out => c207);
	adder0208: full_adder port map(a => p12(7), b => p13(6), c_in => p11(8), s => s208, c_out => c208);
	adder0209: full_adder port map(a => c207, b => c206, c_in => c208, s => s209, c_out => c209);
	adder0210: full_adder port map(a => c204, b => c203, c_in => c205, s => s210, c_out => c210);
	adder0211: full_adder port map(a => p5(15), b => p6(14), c_in => p4(16), s => s211, c_out => c211);
	adder0212: full_adder port map(a => p8(12), b => p9(11), c_in => p7(13), s => s212, c_out => c212);
	adder0213: full_adder port map(a => p11(9), b => p12(8), c_in => p10(10), s => s213, c_out => c213);
	adder0214: full_adder port map(a => p14(6), b => p15(5), c_in => p13(7), s => s214, c_out => c214);
	adder0215: full_adder port map(a => c213, b => c212, c_in => c214, s => s215, c_out => c215);
	adder0216: full_adder port map(a => c210, b => c209, c_in => c211, s => s216, c_out => c216);
	adder0217: full_adder port map(a => p7(14), b => p8(13), c_in => p6(15), s => s217, c_out => c217);
	adder0218: full_adder port map(a => p10(11), b => p11(10), c_in => p9(12), s => s218, c_out => c218);
	adder0219: full_adder port map(a => p13(8), b => p14(7), c_in => p12(9), s => s219, c_out => c219);
	adder0220: full_adder port map(a => p16(5), b => p17(4), c_in => p15(6), s => s220, c_out => c220);
	adder0221: full_adder port map(a => c219, b => c218, c_in => c220, s => s221, c_out => c221);
	adder0222: full_adder port map(a => c216, b => c215, c_in => c217, s => s222, c_out => c222);
	adder0223: full_adder port map(a => p9(13), b => p10(12), c_in => p8(14), s => s223, c_out => c223);
	adder0224: full_adder port map(a => p12(10), b => p13(9), c_in => p11(11), s => s224, c_out => c224);
	adder0225: full_adder port map(a => p15(7), b => p16(6), c_in => p14(8), s => s225, c_out => c225);
	adder0226: full_adder port map(a => p18(4), b => p19(3), c_in => p17(5), s => s226, c_out => c226);
	adder0227: full_adder port map(a => c225, b => c224, c_in => c226, s => s227, c_out => c227);
	adder0228: full_adder port map(a => c222, b => c221, c_in => c223, s => s228, c_out => c228);
	adder0229: full_adder port map(a => p11(12), b => p12(11), c_in => p10(13), s => s229, c_out => c229);
	adder0230: full_adder port map(a => p14(9), b => p15(8), c_in => p13(10), s => s230, c_out => c230);
	adder0231: full_adder port map(a => p17(6), b => p18(5), c_in => p16(7), s => s231, c_out => c231);
	adder0232: full_adder port map(a => p20(3), b => p21(2), c_in => p19(4), s => s232, c_out => c232);
	adder0233: full_adder port map(a => c231, b => c230, c_in => c232, s => s233, c_out => c233);
	adder0234: full_adder port map(a => c228, b => c227, c_in => c229, s => s234, c_out => c234);
	adder0235: full_adder port map(a => p13(11), b => p14(10), c_in => p12(12), s => s235, c_out => c235);
	adder0236: full_adder port map(a => p16(8), b => p17(7), c_in => p15(9), s => s236, c_out => c236);
	adder0237: full_adder port map(a => p19(5), b => p20(4), c_in => p18(6), s => s237, c_out => c237);
	adder0238: full_adder port map(a => p22(2), b => p23(1), c_in => p21(3), s => s238, c_out => c238);
	adder0239: full_adder port map(a => c237, b => c236, c_in => c238, s => s239, c_out => c239);
	adder0240: full_adder port map(a => c234, b => c233, c_in => c235, s => s240, c_out => c240);
	adder0241: full_adder port map(a => p15(10), b => p16(9), c_in => p14(11), s => s241, c_out => c241);
	adder0242: full_adder port map(a => p18(7), b => p19(6), c_in => p17(8), s => s242, c_out => c242);
	adder0243: full_adder port map(a => p21(4), b => p22(3), c_in => p20(5), s => s243, c_out => c243);
	adder0244: full_adder port map(a => p24(1), b => p25(0), c_in => p23(2), s => s244, c_out => c244);
	adder0245: full_adder port map(a => c243, b => c242, c_in => c244, s => s245, c_out => c245);
	adder0246: full_adder port map(a => c240, b => c239, c_in => c241, s => s246, c_out => c246);
	adder0247: full_adder port map(a => p17(9), b => p18(8), c_in => p16(10), s => s247, c_out => c247);
	adder0248: full_adder port map(a => p20(6), b => p21(5), c_in => p19(7), s => s248, c_out => c248);
	adder0249: full_adder port map(a => p23(3), b => p24(2), c_in => p22(4), s => s249, c_out => c249);
	adder0250: full_adder port map(a => p26(0), b => s48, c_in => p25(1), s => s250, c_out => c250);
	adder0251: full_adder port map(a => c249, b => c248, c_in => c250, s => s251, c_out => c251);
	adder0252: full_adder port map(a => c246, b => c245, c_in => c247, s => s252, c_out => c252);
	adder0253: full_adder port map(a => p19(8), b => p20(7), c_in => p18(9), s => s253, c_out => c253);
	adder0254: full_adder port map(a => p22(5), b => p23(4), c_in => p21(6), s => s254, c_out => c254);
	adder0255: full_adder port map(a => p25(2), b => p26(1), c_in => p24(3), s => s255, c_out => c255);
	adder0256: full_adder port map(a => s56, b => s57, c_in => p27(0), s => s256, c_out => c256);
	adder0257: full_adder port map(a => c255, b => c254, c_in => c256, s => s257, c_out => c257);
	adder0258: full_adder port map(a => c252, b => c251, c_in => c253, s => s258, c_out => c258);
	adder0259: full_adder port map(a => p21(7), b => p22(6), c_in => p20(8), s => s259, c_out => c259);
	adder0260: full_adder port map(a => p24(4), b => p25(3), c_in => p23(5), s => s260, c_out => c260);
	adder0261: full_adder port map(a => p27(1), b => p28(0), c_in => p26(2), s => s261, c_out => c261);
	adder0262: full_adder port map(a => s65, b => s66, c_in => s0, s => s262, c_out => c262);
	adder0263: full_adder port map(a => c261, b => c260, c_in => c262, s => s263, c_out => c263);
	adder0264: full_adder port map(a => c258, b => c257, c_in => c259, s => s264, c_out => c264);
	adder0265: full_adder port map(a => p23(6), b => p24(5), c_in => p22(7), s => s265, c_out => c265);
	adder0266: full_adder port map(a => p26(3), b => p27(2), c_in => p25(4), s => s266, c_out => c266);
	adder0267: full_adder port map(a => p29(0), b => s1, c_in => p28(1), s => s267, c_out => c267);
	adder0268: full_adder port map(a => s74, b => s75, c_in => s2, s => s268, c_out => c268);
	adder0269: full_adder port map(a => c267, b => c266, c_in => c268, s => s269, c_out => c269);
	adder0270: full_adder port map(a => c264, b => c263, c_in => c265, s => s270, c_out => c270);
	adder0271: full_adder port map(a => p25(5), b => p26(4), c_in => p24(6), s => s271, c_out => c271);
	adder0272: full_adder port map(a => p28(2), b => p29(1), c_in => p27(3), s => s272, c_out => c272);
	adder0273: full_adder port map(a => s3, b => s4, c_in => p30(0), s => s273, c_out => c273);
	adder0274: full_adder port map(a => s83, b => s84, c_in => s5, s => s274, c_out => c274);
	adder0275: full_adder port map(a => c273, b => c272, c_in => c274, s => s275, c_out => c275);
	adder0276: full_adder port map(a => c270, b => c269, c_in => c271, s => s276, c_out => c276);
	adder0277: full_adder port map(a => p27(4), b => p28(3), c_in => p26(5), s => s277, c_out => c277);
	adder0278: full_adder port map(a => p30(1), b => p31(0), c_in => p29(2), s => s278, c_out => c278);
	adder0279: full_adder port map(a => s7, b => s8, c_in => s6, s => s279, c_out => c279);
	adder0280: full_adder port map(a => s92, b => s93, c_in => s9, s => s280, c_out => c280);
	adder0281: full_adder port map(a => c279, b => c278, c_in => c280, s => s281, c_out => c281);
	adder0282: full_adder port map(a => c276, b => c275, c_in => c277, s => s282, c_out => c282);
	adder0283: full_adder port map(a => p27(5), b => p28(4), c_in => p26(6), s => s283, c_out => c283);
	adder0284: full_adder port map(a => p30(2), b => p31(1), c_in => p29(3), s => s284, c_out => c284);
	adder0285: full_adder port map(a => s11, b => s12, c_in => s10, s => s285, c_out => c285);
	adder0286: full_adder port map(a => s101, b => s102, c_in => s13, s => s286, c_out => c286);
	adder0287: full_adder port map(a => c285, b => c284, c_in => c286, s => s287, c_out => c287);
	adder0288: full_adder port map(a => c282, b => c281, c_in => c283, s => s288, c_out => c288);
	adder0289: full_adder port map(a => p26(7), b => p27(6), c_in => p25(8), s => s289, c_out => c289);
	adder0290: full_adder port map(a => p29(4), b => p30(3), c_in => p28(5), s => s290, c_out => c290);
	adder0291: full_adder port map(a => s14, b => s15, c_in => p31(2), s => s291, c_out => c291);
	adder0292: full_adder port map(a => s110, b => s111, c_in => s16, s => s292, c_out => c292);
	adder0293: full_adder port map(a => c291, b => c290, c_in => c292, s => s293, c_out => c293);
	adder0294: full_adder port map(a => c288, b => c287, c_in => c289, s => s294, c_out => c294);
	adder0295: full_adder port map(a => p25(9), b => p26(8), c_in => p24(10), s => s295, c_out => c295);
	adder0296: full_adder port map(a => p28(6), b => p29(5), c_in => p27(7), s => s296, c_out => c296);
	adder0297: full_adder port map(a => p31(3), b => s17, c_in => p30(4), s => s297, c_out => c297);
	adder0298: full_adder port map(a => s119, b => s120, c_in => s18, s => s298, c_out => c298);
	adder0299: full_adder port map(a => c297, b => c296, c_in => c298, s => s299, c_out => c299);
	adder0300: full_adder port map(a => c294, b => c293, c_in => c295, s => s300, c_out => c300);
	adder0301: full_adder port map(a => p24(11), b => p25(10), c_in => p23(12), s => s301, c_out => c301);
	adder0302: full_adder port map(a => p27(8), b => p28(7), c_in => p26(9), s => s302, c_out => c302);
	adder0303: full_adder port map(a => p30(5), b => p31(4), c_in => p29(6), s => s303, c_out => c303);
	adder0304: full_adder port map(a => s128, b => s129, c_in => s19, s => s304, c_out => c304);
	adder0305: full_adder port map(a => c303, b => c302, c_in => c304, s => s305, c_out => c305);
	adder0306: full_adder port map(a => c300, b => c299, c_in => c301, s => s306, c_out => c306);
	adder0307: full_adder port map(a => p23(13), b => p24(12), c_in => p22(14), s => s307, c_out => c307);
	adder0308: full_adder port map(a => p26(10), b => p27(9), c_in => p25(11), s => s308, c_out => c308);
	adder0309: full_adder port map(a => p29(7), b => p30(6), c_in => p28(8), s => s309, c_out => c309);
	adder0310: full_adder port map(a => s137, b => s138, c_in => p31(5), s => s310, c_out => c310);
	adder0311: full_adder port map(a => c309, b => c308, c_in => c310, s => s311, c_out => c311);
	adder0312: full_adder port map(a => c306, b => c305, c_in => c307, s => s312, c_out => c312);
	adder0313: full_adder port map(a => p22(15), b => p23(14), c_in => p21(16), s => s313, c_out => c313);
	adder0314: full_adder port map(a => p25(12), b => p26(11), c_in => p24(13), s => s314, c_out => c314);
	adder0315: full_adder port map(a => p28(9), b => p29(8), c_in => p27(10), s => s315, c_out => c315);
	adder0316: full_adder port map(a => p31(6), b => s146, c_in => p30(7), s => s316, c_out => c316);
	adder0317: full_adder port map(a => c315, b => c314, c_in => c316, s => s317, c_out => c317);
	adder0318: full_adder port map(a => c312, b => c311, c_in => c313, s => s318, c_out => c318);
	adder0319: full_adder port map(a => p21(17), b => p22(16), c_in => p20(18), s => s319, c_out => c319);
	adder0320: full_adder port map(a => p24(14), b => p25(13), c_in => p23(15), s => s320, c_out => c320);
	adder0321: full_adder port map(a => p27(11), b => p28(10), c_in => p26(12), s => s321, c_out => c321);
	adder0322: full_adder port map(a => p30(8), b => p31(7), c_in => p29(9), s => s322, c_out => c322);
	adder0323: full_adder port map(a => c321, b => c320, c_in => c322, s => s323, c_out => c323);
	adder0324: full_adder port map(a => c318, b => c317, c_in => c319, s => s324, c_out => c324);
	adder0325: full_adder port map(a => p20(19), b => p21(18), c_in => p19(20), s => s325, c_out => c325);
	adder0326: full_adder port map(a => p23(16), b => p24(15), c_in => p22(17), s => s326, c_out => c326);
	adder0327: full_adder port map(a => p26(13), b => p27(12), c_in => p25(14), s => s327, c_out => c327);
	adder0328: full_adder port map(a => p29(10), b => p30(9), c_in => p28(11), s => s328, c_out => c328);
	adder0329: full_adder port map(a => c327, b => c326, c_in => c328, s => s329, c_out => c329);
	adder0330: full_adder port map(a => c324, b => c323, c_in => c325, s => s330, c_out => c330);
	adder0331: full_adder port map(a => p19(21), b => p20(20), c_in => p18(22), s => s331, c_out => c331);
	adder0332: full_adder port map(a => p22(18), b => p23(17), c_in => p21(19), s => s332, c_out => c332);
	adder0333: full_adder port map(a => p25(15), b => p26(14), c_in => p24(16), s => s333, c_out => c333);
	adder0334: full_adder port map(a => p28(12), b => p29(11), c_in => p27(13), s => s334, c_out => c334);
	adder0335: full_adder port map(a => c333, b => c332, c_in => c334, s => s335, c_out => c335);
	adder0336: full_adder port map(a => c330, b => c329, c_in => c331, s => s336, c_out => c336);
	adder0337: full_adder port map(a => p18(23), b => p19(22), c_in => p17(24), s => s337, c_out => c337);
	adder0338: full_adder port map(a => p21(20), b => p22(19), c_in => p20(21), s => s338, c_out => c338);
	adder0339: full_adder port map(a => p24(17), b => p25(16), c_in => p23(18), s => s339, c_out => c339);
	adder0340: full_adder port map(a => p27(14), b => p28(13), c_in => p26(15), s => s340, c_out => c340);
	adder0341: full_adder port map(a => c339, b => c338, c_in => c340, s => s341, c_out => c341);
	adder0342: full_adder port map(a => c336, b => c335, c_in => c337, s => s342, c_out => c342);
	adder0343: full_adder port map(a => p17(25), b => p18(24), c_in => p16(26), s => s343, c_out => c343);
	adder0344: full_adder port map(a => p20(22), b => p21(21), c_in => p19(23), s => s344, c_out => c344);
	adder0345: full_adder port map(a => p23(19), b => p24(18), c_in => p22(20), s => s345, c_out => c345);
	adder0346: full_adder port map(a => p26(16), b => p27(15), c_in => p25(17), s => s346, c_out => c346);
	adder0347: full_adder port map(a => c345, b => c344, c_in => c346, s => s347, c_out => c347);
	adder0348: full_adder port map(a => c342, b => c341, c_in => c343, s => s348, c_out => c348);
	adder0349: full_adder port map(a => p16(27), b => p17(26), c_in => p15(28), s => s349, c_out => c349);
	adder0350: full_adder port map(a => p19(24), b => p20(23), c_in => p18(25), s => s350, c_out => c350);
	adder0351: full_adder port map(a => p22(21), b => p23(20), c_in => p21(22), s => s351, c_out => c351);
	adder0352: full_adder port map(a => p25(18), b => p26(17), c_in => p24(19), s => s352, c_out => c352);
	adder0353: full_adder port map(a => c351, b => c350, c_in => c352, s => s353, c_out => c353);
	adder0354: full_adder port map(a => c348, b => c347, c_in => c349, s => s354, c_out => c354);
	adder0355: full_adder port map(a => p15(29), b => p16(28), c_in => p14(30), s => s355, c_out => c355);
	adder0356: full_adder port map(a => p18(26), b => p19(25), c_in => p17(27), s => s356, c_out => c356);
	adder0357: full_adder port map(a => p21(23), b => p22(22), c_in => p20(24), s => s357, c_out => c357);
	adder0358: full_adder port map(a => p24(20), b => p25(19), c_in => p23(21), s => s358, c_out => c358);
	adder0359: full_adder port map(a => c357, b => c356, c_in => c358, s => s359, c_out => c359);
	adder0360: full_adder port map(a => c354, b => c353, c_in => c355, s => s360, c_out => c360);
	adder0361: full_adder port map(a => p14(31), b => p15(30), c_in => c181, s => s361, c_out => c361);
	adder0362: full_adder port map(a => p17(28), b => p18(27), c_in => p16(29), s => s362, c_out => c362);
	adder0363: full_adder port map(a => p20(25), b => p21(24), c_in => p19(26), s => s363, c_out => c363);
	adder0364: full_adder port map(a => p23(22), b => p24(21), c_in => p22(23), s => s364, c_out => c364);
	adder0365: full_adder port map(a => c363, b => c362, c_in => c364, s => s365, c_out => c365);
	adder0366: full_adder port map(a => c360, b => c359, c_in => c361, s => s366, c_out => c366);
	adder0367: full_adder port map(a => p16(30), b => p17(29), c_in => p15(31), s => s367, c_out => c367);
	adder0368: full_adder port map(a => p19(27), b => p20(26), c_in => p18(28), s => s368, c_out => c368);
	adder0369: full_adder port map(a => p22(24), b => p23(23), c_in => p21(25), s => s369, c_out => c369);
	adder0370: full_adder port map(a => c368, b => c367, c_in => c369, s => s370, c_out => c370);
	adder0371: full_adder port map(a => c365, b => p16(31), c_in => c366, s => s371, c_out => c371);
	adder0372: full_adder port map(a => p18(29), b => p19(28), c_in => p17(30), s => s372, c_out => c372);
	adder0373: full_adder port map(a => p21(26), b => p22(25), c_in => p20(27), s => s373, c_out => c373);
	adder0374: full_adder port map(a => c372, b => c371, c_in => c373, s => s374, c_out => c374);
	adder0375: full_adder port map(a => p17(31), b => p18(30), c_in => c370, s => s375, c_out => c375);
	adder0376: full_adder port map(a => p20(28), b => p21(27), c_in => p19(29), s => s376, c_out => c376);
	adder0377: full_adder port map(a => c375, b => c374, c_in => c376, s => s377, c_out => c377);
	adder0378: full_adder port map(a => p19(30), b => p20(29), c_in => p18(31), s => s378, c_out => c378);
	adder0379: full_adder port map(a => c377, b => p19(31), c_in => c378, s => s379, c_out => c379);
	adder0380: half_adder port map(a => p0(9), b => p1(8), s => s380, c_out => c380);
	adder0381: full_adder port map(a => p0(10), b => p1(9), c_in => c380, s => s381, c_out => c381);
	adder0382: half_adder port map(a => p2(8), b => p3(7), s => s382, c_out => c382);
	adder0383: full_adder port map(a => c381, b => p0(11), c_in => c382, s => s383, c_out => c383);
	adder0384: full_adder port map(a => p2(9), b => p3(8), c_in => p1(10), s => s384, c_out => c384);
	adder0385: half_adder port map(a => p4(7), b => p5(6), s => s385, c_out => c385);
	adder0386: full_adder port map(a => c384, b => c383, c_in => c385, s => s386, c_out => c386);
	adder0387: full_adder port map(a => p1(11), b => p2(10), c_in => p0(12), s => s387, c_out => c387);
	adder0388: full_adder port map(a => p4(8), b => p5(7), c_in => p3(9), s => s388, c_out => c388);
	adder0389: half_adder port map(a => p6(6), b => p7(5), s => s389, c_out => c389);
	adder0390: full_adder port map(a => c388, b => c387, c_in => c389, s => s390, c_out => c390);
	adder0391: full_adder port map(a => p2(11), b => p3(10), c_in => c386, s => s391, c_out => c391);
	adder0392: full_adder port map(a => p5(8), b => p6(7), c_in => p4(9), s => s392, c_out => c392);
	adder0393: full_adder port map(a => p8(5), b => p9(4), c_in => p7(6), s => s393, c_out => c393);
	adder0394: full_adder port map(a => c392, b => c391, c_in => c393, s => s394, c_out => c394);
	adder0395: full_adder port map(a => p4(10), b => p5(9), c_in => c390, s => s395, c_out => c395);
	adder0396: full_adder port map(a => p7(7), b => p8(6), c_in => p6(8), s => s396, c_out => c396);
	adder0397: full_adder port map(a => p10(4), b => p11(3), c_in => p9(5), s => s397, c_out => c397);
	adder0398: full_adder port map(a => c396, b => c395, c_in => c397, s => s398, c_out => c398);
	adder0399: full_adder port map(a => p6(9), b => p7(8), c_in => c394, s => s399, c_out => c399);
	adder0400: full_adder port map(a => p9(6), b => p10(5), c_in => p8(7), s => s400, c_out => c400);
	adder0401: full_adder port map(a => p12(3), b => p13(2), c_in => p11(4), s => s401, c_out => c401);
	adder0402: full_adder port map(a => c400, b => c399, c_in => c401, s => s402, c_out => c402);
	adder0403: full_adder port map(a => p8(8), b => p9(7), c_in => c398, s => s403, c_out => c403);
	adder0404: full_adder port map(a => p11(5), b => p12(4), c_in => p10(6), s => s404, c_out => c404);
	adder0405: full_adder port map(a => p14(2), b => p15(1), c_in => p13(3), s => s405, c_out => c405);
	adder0406: full_adder port map(a => c404, b => c403, c_in => c405, s => s406, c_out => c406);
	adder0407: full_adder port map(a => p10(7), b => p11(6), c_in => c402, s => s407, c_out => c407);
	adder0408: full_adder port map(a => p13(4), b => p14(3), c_in => p12(5), s => s408, c_out => c408);
	adder0409: full_adder port map(a => p16(1), b => p17(0), c_in => p15(2), s => s409, c_out => c409);
	adder0410: full_adder port map(a => c408, b => c407, c_in => c409, s => s410, c_out => c410);
	adder0411: full_adder port map(a => p12(6), b => p13(5), c_in => c406, s => s411, c_out => c411);
	adder0412: full_adder port map(a => p15(3), b => p16(2), c_in => p14(4), s => s412, c_out => c412);
	adder0413: full_adder port map(a => p18(0), b => s197, c_in => p17(1), s => s413, c_out => c413);
	adder0414: full_adder port map(a => c412, b => c411, c_in => c413, s => s414, c_out => c414);
	adder0415: full_adder port map(a => p14(5), b => p15(4), c_in => c410, s => s415, c_out => c415);
	adder0416: full_adder port map(a => p17(2), b => p18(1), c_in => p16(3), s => s416, c_out => c416);
	adder0417: full_adder port map(a => s20, b => s203, c_in => p19(0), s => s417, c_out => c417);
	adder0418: full_adder port map(a => c416, b => c415, c_in => c417, s => s418, c_out => c418);
	adder0419: full_adder port map(a => p16(4), b => p17(3), c_in => c414, s => s419, c_out => c419);
	adder0420: full_adder port map(a => p19(1), b => p20(0), c_in => p18(2), s => s420, c_out => c420);
	adder0421: full_adder port map(a => s22, b => s209, c_in => s21, s => s421, c_out => c421);
	adder0422: full_adder port map(a => c420, b => c419, c_in => c421, s => s422, c_out => c422);
	adder0423: full_adder port map(a => p18(3), b => p19(2), c_in => c418, s => s423, c_out => c423);
	adder0424: full_adder port map(a => p21(0), b => s23, c_in => p20(1), s => s424, c_out => c424);
	adder0425: full_adder port map(a => s25, b => s215, c_in => s24, s => s425, c_out => c425);
	adder0426: full_adder port map(a => c424, b => c423, c_in => c425, s => s426, c_out => c426);
	adder0427: full_adder port map(a => p20(2), b => p21(1), c_in => c422, s => s427, c_out => c427);
	adder0428: full_adder port map(a => s26, b => s27, c_in => p22(0), s => s428, c_out => c428);
	adder0429: full_adder port map(a => s29, b => s221, c_in => s28, s => s429, c_out => c429);
	adder0430: full_adder port map(a => c428, b => c427, c_in => c429, s => s430, c_out => c430);
	adder0431: full_adder port map(a => p22(1), b => p23(0), c_in => c426, s => s431, c_out => c431);
	adder0432: full_adder port map(a => s31, b => s32, c_in => s30, s => s432, c_out => c432);
	adder0433: full_adder port map(a => s34, b => s227, c_in => s33, s => s433, c_out => c433);
	adder0434: full_adder port map(a => c432, b => c431, c_in => c433, s => s434, c_out => c434);
	adder0435: full_adder port map(a => p24(0), b => s35, c_in => c430, s => s435, c_out => c435);
	adder0436: full_adder port map(a => s37, b => s38, c_in => s36, s => s436, c_out => c436);
	adder0437: full_adder port map(a => s40, b => s233, c_in => s39, s => s437, c_out => c437);
	adder0438: full_adder port map(a => c436, b => c435, c_in => c437, s => s438, c_out => c438);
	adder0439: full_adder port map(a => s41, b => s42, c_in => c434, s => s439, c_out => c439);
	adder0440: full_adder port map(a => s44, b => s45, c_in => s43, s => s440, c_out => c440);
	adder0441: full_adder port map(a => s47, b => s239, c_in => s46, s => s441, c_out => c441);
	adder0442: full_adder port map(a => c440, b => c439, c_in => c441, s => s442, c_out => c442);
	adder0443: full_adder port map(a => s49, b => s50, c_in => c438, s => s443, c_out => c443);
	adder0444: full_adder port map(a => s52, b => s53, c_in => s51, s => s444, c_out => c444);
	adder0445: full_adder port map(a => s55, b => s245, c_in => s54, s => s445, c_out => c445);
	adder0446: full_adder port map(a => c444, b => c443, c_in => c445, s => s446, c_out => c446);
	adder0447: full_adder port map(a => s58, b => s59, c_in => c442, s => s447, c_out => c447);
	adder0448: full_adder port map(a => s61, b => s62, c_in => s60, s => s448, c_out => c448);
	adder0449: full_adder port map(a => s64, b => s251, c_in => s63, s => s449, c_out => c449);
	adder0450: full_adder port map(a => c448, b => c447, c_in => c449, s => s450, c_out => c450);
	adder0451: full_adder port map(a => s67, b => s68, c_in => c446, s => s451, c_out => c451);
	adder0452: full_adder port map(a => s70, b => s71, c_in => s69, s => s452, c_out => c452);
	adder0453: full_adder port map(a => s73, b => s257, c_in => s72, s => s453, c_out => c453);
	adder0454: full_adder port map(a => c452, b => c451, c_in => c453, s => s454, c_out => c454);
	adder0455: full_adder port map(a => s76, b => s77, c_in => c450, s => s455, c_out => c455);
	adder0456: full_adder port map(a => s79, b => s80, c_in => s78, s => s456, c_out => c456);
	adder0457: full_adder port map(a => s82, b => s263, c_in => s81, s => s457, c_out => c457);
	adder0458: full_adder port map(a => c456, b => c455, c_in => c457, s => s458, c_out => c458);
	adder0459: full_adder port map(a => s85, b => s86, c_in => c454, s => s459, c_out => c459);
	adder0460: full_adder port map(a => s88, b => s89, c_in => s87, s => s460, c_out => c460);
	adder0461: full_adder port map(a => s91, b => s269, c_in => s90, s => s461, c_out => c461);
	adder0462: full_adder port map(a => c460, b => c459, c_in => c461, s => s462, c_out => c462);
	adder0463: full_adder port map(a => s94, b => s95, c_in => c458, s => s463, c_out => c463);
	adder0464: full_adder port map(a => s97, b => s98, c_in => s96, s => s464, c_out => c464);
	adder0465: full_adder port map(a => s100, b => s275, c_in => s99, s => s465, c_out => c465);
	adder0466: full_adder port map(a => c464, b => c463, c_in => c465, s => s466, c_out => c466);
	adder0467: full_adder port map(a => s103, b => s104, c_in => c462, s => s467, c_out => c467);
	adder0468: full_adder port map(a => s106, b => s107, c_in => s105, s => s468, c_out => c468);
	adder0469: full_adder port map(a => s109, b => s281, c_in => s108, s => s469, c_out => c469);
	adder0470: full_adder port map(a => c468, b => c467, c_in => c469, s => s470, c_out => c470);
	adder0471: full_adder port map(a => s112, b => s113, c_in => c466, s => s471, c_out => c471);
	adder0472: full_adder port map(a => s115, b => s116, c_in => s114, s => s472, c_out => c472);
	adder0473: full_adder port map(a => s118, b => s287, c_in => s117, s => s473, c_out => c473);
	adder0474: full_adder port map(a => c472, b => c471, c_in => c473, s => s474, c_out => c474);
	adder0475: full_adder port map(a => s121, b => s122, c_in => c470, s => s475, c_out => c475);
	adder0476: full_adder port map(a => s124, b => s125, c_in => s123, s => s476, c_out => c476);
	adder0477: full_adder port map(a => s127, b => s293, c_in => s126, s => s477, c_out => c477);
	adder0478: full_adder port map(a => c476, b => c475, c_in => c477, s => s478, c_out => c478);
	adder0479: full_adder port map(a => s130, b => s131, c_in => c474, s => s479, c_out => c479);
	adder0480: full_adder port map(a => s133, b => s134, c_in => s132, s => s480, c_out => c480);
	adder0481: full_adder port map(a => s136, b => s299, c_in => s135, s => s481, c_out => c481);
	adder0482: full_adder port map(a => c480, b => c479, c_in => c481, s => s482, c_out => c482);
	adder0483: full_adder port map(a => s139, b => s140, c_in => c478, s => s483, c_out => c483);
	adder0484: full_adder port map(a => s142, b => s143, c_in => s141, s => s484, c_out => c484);
	adder0485: full_adder port map(a => s145, b => s305, c_in => s144, s => s485, c_out => c485);
	adder0486: full_adder port map(a => c484, b => c483, c_in => c485, s => s486, c_out => c486);
	adder0487: full_adder port map(a => s147, b => s148, c_in => c482, s => s487, c_out => c487);
	adder0488: full_adder port map(a => s150, b => s151, c_in => s149, s => s488, c_out => c488);
	adder0489: full_adder port map(a => s153, b => s311, c_in => s152, s => s489, c_out => c489);
	adder0490: full_adder port map(a => c488, b => c487, c_in => c489, s => s490, c_out => c490);
	adder0491: full_adder port map(a => s154, b => s155, c_in => c486, s => s491, c_out => c491);
	adder0492: full_adder port map(a => s157, b => s158, c_in => s156, s => s492, c_out => c492);
	adder0493: full_adder port map(a => s160, b => s317, c_in => s159, s => s493, c_out => c493);
	adder0494: full_adder port map(a => c492, b => c491, c_in => c493, s => s494, c_out => c494);
	adder0495: full_adder port map(a => p31(8), b => s161, c_in => c490, s => s495, c_out => c495);
	adder0496: full_adder port map(a => s163, b => s164, c_in => s162, s => s496, c_out => c496);
	adder0497: full_adder port map(a => s166, b => s323, c_in => s165, s => s497, c_out => c497);
	adder0498: full_adder port map(a => c496, b => c495, c_in => c497, s => s498, c_out => c498);
	adder0499: full_adder port map(a => p30(10), b => p31(9), c_in => c494, s => s499, c_out => c499);
	adder0500: full_adder port map(a => s168, b => s169, c_in => s167, s => s500, c_out => c500);
	adder0501: full_adder port map(a => s171, b => s329, c_in => s170, s => s501, c_out => c501);
	adder0502: full_adder port map(a => c500, b => c499, c_in => c501, s => s502, c_out => c502);
	adder0503: full_adder port map(a => p29(12), b => p30(11), c_in => c498, s => s503, c_out => c503);
	adder0504: full_adder port map(a => s172, b => s173, c_in => p31(10), s => s504, c_out => c504);
	adder0505: full_adder port map(a => s175, b => s335, c_in => s174, s => s505, c_out => c505);
	adder0506: full_adder port map(a => c504, b => c503, c_in => c505, s => s506, c_out => c506);
	adder0507: full_adder port map(a => p28(14), b => p29(13), c_in => c502, s => s507, c_out => c507);
	adder0508: full_adder port map(a => p31(11), b => s176, c_in => p30(12), s => s508, c_out => c508);
	adder0509: full_adder port map(a => s178, b => s341, c_in => s177, s => s509, c_out => c509);
	adder0510: full_adder port map(a => c508, b => c507, c_in => c509, s => s510, c_out => c510);
	adder0511: full_adder port map(a => p27(16), b => p28(15), c_in => c506, s => s511, c_out => c511);
	adder0512: full_adder port map(a => p30(13), b => p31(12), c_in => p29(14), s => s512, c_out => c512);
	adder0513: full_adder port map(a => s180, b => s347, c_in => s179, s => s513, c_out => c513);
	adder0514: full_adder port map(a => c512, b => c511, c_in => c513, s => s514, c_out => c514);
	adder0515: full_adder port map(a => p26(18), b => p27(17), c_in => c510, s => s515, c_out => c515);
	adder0516: full_adder port map(a => p29(15), b => p30(14), c_in => p28(16), s => s516, c_out => c516);
	adder0517: full_adder port map(a => s181, b => s353, c_in => p31(13), s => s517, c_out => c517);
	adder0518: full_adder port map(a => c516, b => c515, c_in => c517, s => s518, c_out => c518);
	adder0519: full_adder port map(a => p25(20), b => p26(19), c_in => c514, s => s519, c_out => c519);
	adder0520: full_adder port map(a => p28(17), b => p29(16), c_in => p27(18), s => s520, c_out => c520);
	adder0521: full_adder port map(a => p31(14), b => s359, c_in => p30(15), s => s521, c_out => c521);
	adder0522: full_adder port map(a => c520, b => c519, c_in => c521, s => s522, c_out => c522);
	adder0523: full_adder port map(a => p24(22), b => p25(21), c_in => c518, s => s523, c_out => c523);
	adder0524: full_adder port map(a => p27(19), b => p28(18), c_in => p26(20), s => s524, c_out => c524);
	adder0525: full_adder port map(a => p30(16), b => p31(15), c_in => p29(17), s => s525, c_out => c525);
	adder0526: full_adder port map(a => c524, b => c523, c_in => c525, s => s526, c_out => c526);
	adder0527: full_adder port map(a => p23(24), b => p24(23), c_in => c522, s => s527, c_out => c527);
	adder0528: full_adder port map(a => p26(21), b => p27(20), c_in => p25(22), s => s528, c_out => c528);
	adder0529: full_adder port map(a => p29(18), b => p30(17), c_in => p28(19), s => s529, c_out => c529);
	adder0530: full_adder port map(a => c528, b => c527, c_in => c529, s => s530, c_out => c530);
	adder0531: full_adder port map(a => p22(26), b => p23(25), c_in => c526, s => s531, c_out => c531);
	adder0532: full_adder port map(a => p25(23), b => p26(22), c_in => p24(24), s => s532, c_out => c532);
	adder0533: full_adder port map(a => p28(20), b => p29(19), c_in => p27(21), s => s533, c_out => c533);
	adder0534: full_adder port map(a => c532, b => c531, c_in => c533, s => s534, c_out => c534);
	adder0535: full_adder port map(a => p21(28), b => p22(27), c_in => c530, s => s535, c_out => c535);
	adder0536: full_adder port map(a => p24(25), b => p25(24), c_in => p23(26), s => s536, c_out => c536);
	adder0537: full_adder port map(a => p27(22), b => p28(21), c_in => p26(23), s => s537, c_out => c537);
	adder0538: full_adder port map(a => c536, b => c535, c_in => c537, s => s538, c_out => c538);
	adder0539: full_adder port map(a => p20(30), b => p21(29), c_in => c534, s => s539, c_out => c539);
	adder0540: full_adder port map(a => p23(27), b => p24(26), c_in => p22(28), s => s540, c_out => c540);
	adder0541: full_adder port map(a => p26(24), b => p27(23), c_in => p25(25), s => s541, c_out => c541);
	adder0542: full_adder port map(a => c540, b => c539, c_in => c541, s => s542, c_out => c542);
	adder0543: full_adder port map(a => c379, b => p20(31), c_in => c538, s => s543, c_out => c543);
	adder0544: full_adder port map(a => p22(29), b => p23(28), c_in => p21(30), s => s544, c_out => c544);
	adder0545: full_adder port map(a => p25(26), b => p26(25), c_in => p24(27), s => s545, c_out => c545);
	adder0546: full_adder port map(a => c544, b => c543, c_in => c545, s => s546, c_out => c546);
	adder0547: full_adder port map(a => p21(31), b => p22(30), c_in => c542, s => s547, c_out => c547);
	adder0548: full_adder port map(a => p24(28), b => p25(27), c_in => p23(29), s => s548, c_out => c548);
	adder0549: full_adder port map(a => c547, b => c546, c_in => c548, s => s549, c_out => c549);
	adder0550: full_adder port map(a => p23(30), b => p24(29), c_in => p22(31), s => s550, c_out => c550);
	adder0551: full_adder port map(a => c549, b => p23(31), c_in => c550, s => s551, c_out => c551);
	adder0552: half_adder port map(a => p0(6), b => p1(5), s => s552, c_out => c552);
	adder0553: full_adder port map(a => p0(7), b => p1(6), c_in => c552, s => s553, c_out => c553);
	adder0554: half_adder port map(a => p2(5), b => p3(4), s => s554, c_out => c554);
	adder0555: full_adder port map(a => c553, b => p0(8), c_in => c554, s => s555, c_out => c555);
	adder0556: full_adder port map(a => p2(6), b => p3(5), c_in => p1(7), s => s556, c_out => c556);
	adder0557: half_adder port map(a => p4(4), b => p5(3), s => s557, c_out => c557);
	adder0558: full_adder port map(a => c556, b => c555, c_in => c557, s => s558, c_out => c558);
	adder0559: full_adder port map(a => p3(6), b => p4(5), c_in => p2(7), s => s559, c_out => c559);
	adder0560: full_adder port map(a => p6(3), b => p7(2), c_in => p5(4), s => s560, c_out => c560);
	adder0561: full_adder port map(a => c559, b => c558, c_in => c560, s => s561, c_out => c561);
	adder0562: full_adder port map(a => p5(5), b => p6(4), c_in => p4(6), s => s562, c_out => c562);
	adder0563: full_adder port map(a => p8(2), b => p9(1), c_in => p7(3), s => s563, c_out => c563);
	adder0564: full_adder port map(a => c562, b => c561, c_in => c563, s => s564, c_out => c564);
	adder0565: full_adder port map(a => p7(4), b => p8(3), c_in => p6(5), s => s565, c_out => c565);
	adder0566: full_adder port map(a => p10(1), b => p11(0), c_in => p9(2), s => s566, c_out => c566);
	adder0567: full_adder port map(a => c565, b => c564, c_in => c566, s => s567, c_out => c567);
	adder0568: full_adder port map(a => p9(3), b => p10(2), c_in => p8(4), s => s568, c_out => c568);
	adder0569: full_adder port map(a => p12(0), b => s386, c_in => p11(1), s => s569, c_out => c569);
	adder0570: full_adder port map(a => c568, b => c567, c_in => c569, s => s570, c_out => c570);
	adder0571: full_adder port map(a => p11(2), b => p12(1), c_in => p10(3), s => s571, c_out => c571);
	adder0572: full_adder port map(a => s182, b => s390, c_in => p13(0), s => s572, c_out => c572);
	adder0573: full_adder port map(a => c571, b => c570, c_in => c572, s => s573, c_out => c573);
	adder0574: full_adder port map(a => p13(1), b => p14(0), c_in => p12(2), s => s574, c_out => c574);
	adder0575: full_adder port map(a => s184, b => s394, c_in => s183, s => s575, c_out => c575);
	adder0576: full_adder port map(a => c574, b => c573, c_in => c575, s => s576, c_out => c576);
	adder0577: full_adder port map(a => p15(0), b => s185, c_in => p14(1), s => s577, c_out => c577);
	adder0578: full_adder port map(a => s187, b => s398, c_in => s186, s => s578, c_out => c578);
	adder0579: full_adder port map(a => c577, b => c576, c_in => c578, s => s579, c_out => c579);
	adder0580: full_adder port map(a => s188, b => s189, c_in => p16(0), s => s580, c_out => c580);
	adder0581: full_adder port map(a => s191, b => s402, c_in => s190, s => s581, c_out => c581);
	adder0582: full_adder port map(a => c580, b => c579, c_in => c581, s => s582, c_out => c582);
	adder0583: full_adder port map(a => s193, b => s194, c_in => s192, s => s583, c_out => c583);
	adder0584: full_adder port map(a => s196, b => s406, c_in => s195, s => s584, c_out => c584);
	adder0585: full_adder port map(a => c583, b => c582, c_in => c584, s => s585, c_out => c585);
	adder0586: full_adder port map(a => s199, b => s200, c_in => s198, s => s586, c_out => c586);
	adder0587: full_adder port map(a => s202, b => s410, c_in => s201, s => s587, c_out => c587);
	adder0588: full_adder port map(a => c586, b => c585, c_in => c587, s => s588, c_out => c588);
	adder0589: full_adder port map(a => s205, b => s206, c_in => s204, s => s589, c_out => c589);
	adder0590: full_adder port map(a => s208, b => s414, c_in => s207, s => s590, c_out => c590);
	adder0591: full_adder port map(a => c589, b => c588, c_in => c590, s => s591, c_out => c591);
	adder0592: full_adder port map(a => s211, b => s212, c_in => s210, s => s592, c_out => c592);
	adder0593: full_adder port map(a => s214, b => s418, c_in => s213, s => s593, c_out => c593);
	adder0594: full_adder port map(a => c592, b => c591, c_in => c593, s => s594, c_out => c594);
	adder0595: full_adder port map(a => s217, b => s218, c_in => s216, s => s595, c_out => c595);
	adder0596: full_adder port map(a => s220, b => s422, c_in => s219, s => s596, c_out => c596);
	adder0597: full_adder port map(a => c595, b => c594, c_in => c596, s => s597, c_out => c597);
	adder0598: full_adder port map(a => s223, b => s224, c_in => s222, s => s598, c_out => c598);
	adder0599: full_adder port map(a => s226, b => s426, c_in => s225, s => s599, c_out => c599);
	adder0600: full_adder port map(a => c598, b => c597, c_in => c599, s => s600, c_out => c600);
	adder0601: full_adder port map(a => s229, b => s230, c_in => s228, s => s601, c_out => c601);
	adder0602: full_adder port map(a => s232, b => s430, c_in => s231, s => s602, c_out => c602);
	adder0603: full_adder port map(a => c601, b => c600, c_in => c602, s => s603, c_out => c603);
	adder0604: full_adder port map(a => s235, b => s236, c_in => s234, s => s604, c_out => c604);
	adder0605: full_adder port map(a => s238, b => s434, c_in => s237, s => s605, c_out => c605);
	adder0606: full_adder port map(a => c604, b => c603, c_in => c605, s => s606, c_out => c606);
	adder0607: full_adder port map(a => s241, b => s242, c_in => s240, s => s607, c_out => c607);
	adder0608: full_adder port map(a => s244, b => s438, c_in => s243, s => s608, c_out => c608);
	adder0609: full_adder port map(a => c607, b => c606, c_in => c608, s => s609, c_out => c609);
	adder0610: full_adder port map(a => s247, b => s248, c_in => s246, s => s610, c_out => c610);
	adder0611: full_adder port map(a => s250, b => s442, c_in => s249, s => s611, c_out => c611);
	adder0612: full_adder port map(a => c610, b => c609, c_in => c611, s => s612, c_out => c612);
	adder0613: full_adder port map(a => s253, b => s254, c_in => s252, s => s613, c_out => c613);
	adder0614: full_adder port map(a => s256, b => s446, c_in => s255, s => s614, c_out => c614);
	adder0615: full_adder port map(a => c613, b => c612, c_in => c614, s => s615, c_out => c615);
	adder0616: full_adder port map(a => s259, b => s260, c_in => s258, s => s616, c_out => c616);
	adder0617: full_adder port map(a => s262, b => s450, c_in => s261, s => s617, c_out => c617);
	adder0618: full_adder port map(a => c616, b => c615, c_in => c617, s => s618, c_out => c618);
	adder0619: full_adder port map(a => s265, b => s266, c_in => s264, s => s619, c_out => c619);
	adder0620: full_adder port map(a => s268, b => s454, c_in => s267, s => s620, c_out => c620);
	adder0621: full_adder port map(a => c619, b => c618, c_in => c620, s => s621, c_out => c621);
	adder0622: full_adder port map(a => s271, b => s272, c_in => s270, s => s622, c_out => c622);
	adder0623: full_adder port map(a => s274, b => s458, c_in => s273, s => s623, c_out => c623);
	adder0624: full_adder port map(a => c622, b => c621, c_in => c623, s => s624, c_out => c624);
	adder0625: full_adder port map(a => s277, b => s278, c_in => s276, s => s625, c_out => c625);
	adder0626: full_adder port map(a => s280, b => s462, c_in => s279, s => s626, c_out => c626);
	adder0627: full_adder port map(a => c625, b => c624, c_in => c626, s => s627, c_out => c627);
	adder0628: full_adder port map(a => s283, b => s284, c_in => s282, s => s628, c_out => c628);
	adder0629: full_adder port map(a => s286, b => s466, c_in => s285, s => s629, c_out => c629);
	adder0630: full_adder port map(a => c628, b => c627, c_in => c629, s => s630, c_out => c630);
	adder0631: full_adder port map(a => s289, b => s290, c_in => s288, s => s631, c_out => c631);
	adder0632: full_adder port map(a => s292, b => s470, c_in => s291, s => s632, c_out => c632);
	adder0633: full_adder port map(a => c631, b => c630, c_in => c632, s => s633, c_out => c633);
	adder0634: full_adder port map(a => s295, b => s296, c_in => s294, s => s634, c_out => c634);
	adder0635: full_adder port map(a => s298, b => s474, c_in => s297, s => s635, c_out => c635);
	adder0636: full_adder port map(a => c634, b => c633, c_in => c635, s => s636, c_out => c636);
	adder0637: full_adder port map(a => s301, b => s302, c_in => s300, s => s637, c_out => c637);
	adder0638: full_adder port map(a => s304, b => s478, c_in => s303, s => s638, c_out => c638);
	adder0639: full_adder port map(a => c637, b => c636, c_in => c638, s => s639, c_out => c639);
	adder0640: full_adder port map(a => s307, b => s308, c_in => s306, s => s640, c_out => c640);
	adder0641: full_adder port map(a => s310, b => s482, c_in => s309, s => s641, c_out => c641);
	adder0642: full_adder port map(a => c640, b => c639, c_in => c641, s => s642, c_out => c642);
	adder0643: full_adder port map(a => s313, b => s314, c_in => s312, s => s643, c_out => c643);
	adder0644: full_adder port map(a => s316, b => s486, c_in => s315, s => s644, c_out => c644);
	adder0645: full_adder port map(a => c643, b => c642, c_in => c644, s => s645, c_out => c645);
	adder0646: full_adder port map(a => s319, b => s320, c_in => s318, s => s646, c_out => c646);
	adder0647: full_adder port map(a => s322, b => s490, c_in => s321, s => s647, c_out => c647);
	adder0648: full_adder port map(a => c646, b => c645, c_in => c647, s => s648, c_out => c648);
	adder0649: full_adder port map(a => s325, b => s326, c_in => s324, s => s649, c_out => c649);
	adder0650: full_adder port map(a => s328, b => s494, c_in => s327, s => s650, c_out => c650);
	adder0651: full_adder port map(a => c649, b => c648, c_in => c650, s => s651, c_out => c651);
	adder0652: full_adder port map(a => s331, b => s332, c_in => s330, s => s652, c_out => c652);
	adder0653: full_adder port map(a => s334, b => s498, c_in => s333, s => s653, c_out => c653);
	adder0654: full_adder port map(a => c652, b => c651, c_in => c653, s => s654, c_out => c654);
	adder0655: full_adder port map(a => s337, b => s338, c_in => s336, s => s655, c_out => c655);
	adder0656: full_adder port map(a => s340, b => s502, c_in => s339, s => s656, c_out => c656);
	adder0657: full_adder port map(a => c655, b => c654, c_in => c656, s => s657, c_out => c657);
	adder0658: full_adder port map(a => s343, b => s344, c_in => s342, s => s658, c_out => c658);
	adder0659: full_adder port map(a => s346, b => s506, c_in => s345, s => s659, c_out => c659);
	adder0660: full_adder port map(a => c658, b => c657, c_in => c659, s => s660, c_out => c660);
	adder0661: full_adder port map(a => s349, b => s350, c_in => s348, s => s661, c_out => c661);
	adder0662: full_adder port map(a => s352, b => s510, c_in => s351, s => s662, c_out => c662);
	adder0663: full_adder port map(a => c661, b => c660, c_in => c662, s => s663, c_out => c663);
	adder0664: full_adder port map(a => s355, b => s356, c_in => s354, s => s664, c_out => c664);
	adder0665: full_adder port map(a => s358, b => s514, c_in => s357, s => s665, c_out => c665);
	adder0666: full_adder port map(a => c664, b => c663, c_in => c665, s => s666, c_out => c666);
	adder0667: full_adder port map(a => s361, b => s362, c_in => s360, s => s667, c_out => c667);
	adder0668: full_adder port map(a => s364, b => s518, c_in => s363, s => s668, c_out => c668);
	adder0669: full_adder port map(a => c667, b => c666, c_in => c668, s => s669, c_out => c669);
	adder0670: full_adder port map(a => s366, b => s367, c_in => s365, s => s670, c_out => c670);
	adder0671: full_adder port map(a => s369, b => s522, c_in => s368, s => s671, c_out => c671);
	adder0672: full_adder port map(a => c670, b => c669, c_in => c671, s => s672, c_out => c672);
	adder0673: full_adder port map(a => s370, b => s371, c_in => p31(16), s => s673, c_out => c673);
	adder0674: full_adder port map(a => s373, b => s526, c_in => s372, s => s674, c_out => c674);
	adder0675: full_adder port map(a => c673, b => c672, c_in => c674, s => s675, c_out => c675);
	adder0676: full_adder port map(a => p31(17), b => s374, c_in => p30(18), s => s676, c_out => c676);
	adder0677: full_adder port map(a => s376, b => s530, c_in => s375, s => s677, c_out => c677);
	adder0678: full_adder port map(a => c676, b => c675, c_in => c677, s => s678, c_out => c678);
	adder0679: full_adder port map(a => p30(19), b => p31(18), c_in => p29(20), s => s679, c_out => c679);
	adder0680: full_adder port map(a => s378, b => s534, c_in => s377, s => s680, c_out => c680);
	adder0681: full_adder port map(a => c679, b => c678, c_in => c680, s => s681, c_out => c681);
	adder0682: full_adder port map(a => p29(21), b => p30(20), c_in => p28(22), s => s682, c_out => c682);
	adder0683: full_adder port map(a => s379, b => s538, c_in => p31(19), s => s683, c_out => c683);
	adder0684: full_adder port map(a => c682, b => c681, c_in => c683, s => s684, c_out => c684);
	adder0685: full_adder port map(a => p28(23), b => p29(22), c_in => p27(24), s => s685, c_out => c685);
	adder0686: full_adder port map(a => p31(20), b => s542, c_in => p30(21), s => s686, c_out => c686);
	adder0687: full_adder port map(a => c685, b => c684, c_in => c686, s => s687, c_out => c687);
	adder0688: full_adder port map(a => p27(25), b => p28(24), c_in => p26(26), s => s688, c_out => c688);
	adder0689: full_adder port map(a => p30(22), b => p31(21), c_in => p29(23), s => s689, c_out => c689);
	adder0690: full_adder port map(a => c688, b => c687, c_in => c689, s => s690, c_out => c690);
	adder0691: full_adder port map(a => p26(27), b => p27(26), c_in => p25(28), s => s691, c_out => c691);
	adder0692: full_adder port map(a => p29(24), b => p30(23), c_in => p28(25), s => s692, c_out => c692);
	adder0693: full_adder port map(a => c691, b => c690, c_in => c692, s => s693, c_out => c693);
	adder0694: full_adder port map(a => p25(29), b => p26(28), c_in => p24(30), s => s694, c_out => c694);
	adder0695: full_adder port map(a => p28(26), b => p29(25), c_in => p27(27), s => s695, c_out => c695);
	adder0696: full_adder port map(a => c694, b => c693, c_in => c695, s => s696, c_out => c696);
	adder0697: full_adder port map(a => p24(31), b => p25(30), c_in => c551, s => s697, c_out => c697);
	adder0698: full_adder port map(a => p27(28), b => p28(27), c_in => p26(29), s => s698, c_out => c698);
	adder0699: full_adder port map(a => c697, b => c696, c_in => c698, s => s699, c_out => c699);
	adder0700: full_adder port map(a => p26(30), b => p27(29), c_in => p25(31), s => s700, c_out => c700);
	adder0701: full_adder port map(a => c699, b => p26(31), c_in => c700, s => s701, c_out => c701);
	adder0702: half_adder port map(a => p0(4), b => p1(3), s => s702, c_out => c702);
	adder0703: full_adder port map(a => p0(5), b => p1(4), c_in => c702, s => s703, c_out => c703);
	adder0704: half_adder port map(a => p2(3), b => p3(2), s => s704, c_out => c704);
	adder0705: full_adder port map(a => c703, b => p2(4), c_in => c704, s => s705, c_out => c705);
	adder0706: full_adder port map(a => p4(2), b => p5(1), c_in => p3(3), s => s706, c_out => c706);
	adder0707: full_adder port map(a => c705, b => p4(3), c_in => c706, s => s707, c_out => c707);
	adder0708: full_adder port map(a => p6(1), b => p7(0), c_in => p5(2), s => s708, c_out => c708);
	adder0709: full_adder port map(a => c707, b => p6(2), c_in => c708, s => s709, c_out => c709);
	adder0710: full_adder port map(a => p8(0), b => s555, c_in => p7(1), s => s710, c_out => c710);
	adder0711: full_adder port map(a => c709, b => p8(1), c_in => c710, s => s711, c_out => c711);
	adder0712: full_adder port map(a => s380, b => s558, c_in => p9(0), s => s712, c_out => c712);
	adder0713: full_adder port map(a => c711, b => p10(0), c_in => c712, s => s713, c_out => c713);
	adder0714: full_adder port map(a => s382, b => s561, c_in => s381, s => s714, c_out => c714);
	adder0715: full_adder port map(a => c713, b => s383, c_in => c714, s => s715, c_out => c715);
	adder0716: full_adder port map(a => s385, b => s564, c_in => s384, s => s716, c_out => c716);
	adder0717: full_adder port map(a => c715, b => s387, c_in => c716, s => s717, c_out => c717);
	adder0718: full_adder port map(a => s389, b => s567, c_in => s388, s => s718, c_out => c718);
	adder0719: full_adder port map(a => c717, b => s391, c_in => c718, s => s719, c_out => c719);
	adder0720: full_adder port map(a => s393, b => s570, c_in => s392, s => s720, c_out => c720);
	adder0721: full_adder port map(a => c719, b => s395, c_in => c720, s => s721, c_out => c721);
	adder0722: full_adder port map(a => s397, b => s573, c_in => s396, s => s722, c_out => c722);
	adder0723: full_adder port map(a => c721, b => s399, c_in => c722, s => s723, c_out => c723);
	adder0724: full_adder port map(a => s401, b => s576, c_in => s400, s => s724, c_out => c724);
	adder0725: full_adder port map(a => c723, b => s403, c_in => c724, s => s725, c_out => c725);
	adder0726: full_adder port map(a => s405, b => s579, c_in => s404, s => s726, c_out => c726);
	adder0727: full_adder port map(a => c725, b => s407, c_in => c726, s => s727, c_out => c727);
	adder0728: full_adder port map(a => s409, b => s582, c_in => s408, s => s728, c_out => c728);
	adder0729: full_adder port map(a => c727, b => s411, c_in => c728, s => s729, c_out => c729);
	adder0730: full_adder port map(a => s413, b => s585, c_in => s412, s => s730, c_out => c730);
	adder0731: full_adder port map(a => c729, b => s415, c_in => c730, s => s731, c_out => c731);
	adder0732: full_adder port map(a => s417, b => s588, c_in => s416, s => s732, c_out => c732);
	adder0733: full_adder port map(a => c731, b => s419, c_in => c732, s => s733, c_out => c733);
	adder0734: full_adder port map(a => s421, b => s591, c_in => s420, s => s734, c_out => c734);
	adder0735: full_adder port map(a => c733, b => s423, c_in => c734, s => s735, c_out => c735);
	adder0736: full_adder port map(a => s425, b => s594, c_in => s424, s => s736, c_out => c736);
	adder0737: full_adder port map(a => c735, b => s427, c_in => c736, s => s737, c_out => c737);
	adder0738: full_adder port map(a => s429, b => s597, c_in => s428, s => s738, c_out => c738);
	adder0739: full_adder port map(a => c737, b => s431, c_in => c738, s => s739, c_out => c739);
	adder0740: full_adder port map(a => s433, b => s600, c_in => s432, s => s740, c_out => c740);
	adder0741: full_adder port map(a => c739, b => s435, c_in => c740, s => s741, c_out => c741);
	adder0742: full_adder port map(a => s437, b => s603, c_in => s436, s => s742, c_out => c742);
	adder0743: full_adder port map(a => c741, b => s439, c_in => c742, s => s743, c_out => c743);
	adder0744: full_adder port map(a => s441, b => s606, c_in => s440, s => s744, c_out => c744);
	adder0745: full_adder port map(a => c743, b => s443, c_in => c744, s => s745, c_out => c745);
	adder0746: full_adder port map(a => s445, b => s609, c_in => s444, s => s746, c_out => c746);
	adder0747: full_adder port map(a => c745, b => s447, c_in => c746, s => s747, c_out => c747);
	adder0748: full_adder port map(a => s449, b => s612, c_in => s448, s => s748, c_out => c748);
	adder0749: full_adder port map(a => c747, b => s451, c_in => c748, s => s749, c_out => c749);
	adder0750: full_adder port map(a => s453, b => s615, c_in => s452, s => s750, c_out => c750);
	adder0751: full_adder port map(a => c749, b => s455, c_in => c750, s => s751, c_out => c751);
	adder0752: full_adder port map(a => s457, b => s618, c_in => s456, s => s752, c_out => c752);
	adder0753: full_adder port map(a => c751, b => s459, c_in => c752, s => s753, c_out => c753);
	adder0754: full_adder port map(a => s461, b => s621, c_in => s460, s => s754, c_out => c754);
	adder0755: full_adder port map(a => c753, b => s463, c_in => c754, s => s755, c_out => c755);
	adder0756: full_adder port map(a => s465, b => s624, c_in => s464, s => s756, c_out => c756);
	adder0757: full_adder port map(a => c755, b => s467, c_in => c756, s => s757, c_out => c757);
	adder0758: full_adder port map(a => s469, b => s627, c_in => s468, s => s758, c_out => c758);
	adder0759: full_adder port map(a => c757, b => s471, c_in => c758, s => s759, c_out => c759);
	adder0760: full_adder port map(a => s473, b => s630, c_in => s472, s => s760, c_out => c760);
	adder0761: full_adder port map(a => c759, b => s475, c_in => c760, s => s761, c_out => c761);
	adder0762: full_adder port map(a => s477, b => s633, c_in => s476, s => s762, c_out => c762);
	adder0763: full_adder port map(a => c761, b => s479, c_in => c762, s => s763, c_out => c763);
	adder0764: full_adder port map(a => s481, b => s636, c_in => s480, s => s764, c_out => c764);
	adder0765: full_adder port map(a => c763, b => s483, c_in => c764, s => s765, c_out => c765);
	adder0766: full_adder port map(a => s485, b => s639, c_in => s484, s => s766, c_out => c766);
	adder0767: full_adder port map(a => c765, b => s487, c_in => c766, s => s767, c_out => c767);
	adder0768: full_adder port map(a => s489, b => s642, c_in => s488, s => s768, c_out => c768);
	adder0769: full_adder port map(a => c767, b => s491, c_in => c768, s => s769, c_out => c769);
	adder0770: full_adder port map(a => s493, b => s645, c_in => s492, s => s770, c_out => c770);
	adder0771: full_adder port map(a => c769, b => s495, c_in => c770, s => s771, c_out => c771);
	adder0772: full_adder port map(a => s497, b => s648, c_in => s496, s => s772, c_out => c772);
	adder0773: full_adder port map(a => c771, b => s499, c_in => c772, s => s773, c_out => c773);
	adder0774: full_adder port map(a => s501, b => s651, c_in => s500, s => s774, c_out => c774);
	adder0775: full_adder port map(a => c773, b => s503, c_in => c774, s => s775, c_out => c775);
	adder0776: full_adder port map(a => s505, b => s654, c_in => s504, s => s776, c_out => c776);
	adder0777: full_adder port map(a => c775, b => s507, c_in => c776, s => s777, c_out => c777);
	adder0778: full_adder port map(a => s509, b => s657, c_in => s508, s => s778, c_out => c778);
	adder0779: full_adder port map(a => c777, b => s511, c_in => c778, s => s779, c_out => c779);
	adder0780: full_adder port map(a => s513, b => s660, c_in => s512, s => s780, c_out => c780);
	adder0781: full_adder port map(a => c779, b => s515, c_in => c780, s => s781, c_out => c781);
	adder0782: full_adder port map(a => s517, b => s663, c_in => s516, s => s782, c_out => c782);
	adder0783: full_adder port map(a => c781, b => s519, c_in => c782, s => s783, c_out => c783);
	adder0784: full_adder port map(a => s521, b => s666, c_in => s520, s => s784, c_out => c784);
	adder0785: full_adder port map(a => c783, b => s523, c_in => c784, s => s785, c_out => c785);
	adder0786: full_adder port map(a => s525, b => s669, c_in => s524, s => s786, c_out => c786);
	adder0787: full_adder port map(a => c785, b => s527, c_in => c786, s => s787, c_out => c787);
	adder0788: full_adder port map(a => s529, b => s672, c_in => s528, s => s788, c_out => c788);
	adder0789: full_adder port map(a => c787, b => s531, c_in => c788, s => s789, c_out => c789);
	adder0790: full_adder port map(a => s533, b => s675, c_in => s532, s => s790, c_out => c790);
	adder0791: full_adder port map(a => c789, b => s535, c_in => c790, s => s791, c_out => c791);
	adder0792: full_adder port map(a => s537, b => s678, c_in => s536, s => s792, c_out => c792);
	adder0793: full_adder port map(a => c791, b => s539, c_in => c792, s => s793, c_out => c793);
	adder0794: full_adder port map(a => s541, b => s681, c_in => s540, s => s794, c_out => c794);
	adder0795: full_adder port map(a => c793, b => s543, c_in => c794, s => s795, c_out => c795);
	adder0796: full_adder port map(a => s545, b => s684, c_in => s544, s => s796, c_out => c796);
	adder0797: full_adder port map(a => c795, b => s546, c_in => c796, s => s797, c_out => c797);
	adder0798: full_adder port map(a => s548, b => s687, c_in => s547, s => s798, c_out => c798);
	adder0799: full_adder port map(a => c797, b => p31(22), c_in => c798, s => s799, c_out => c799);
	adder0800: full_adder port map(a => s550, b => s690, c_in => s549, s => s800, c_out => c800);
	adder0801: full_adder port map(a => c799, b => p30(24), c_in => c800, s => s801, c_out => c801);
	adder0802: full_adder port map(a => s551, b => s693, c_in => p31(23), s => s802, c_out => c802);
	adder0803: full_adder port map(a => c801, b => p29(26), c_in => c802, s => s803, c_out => c803);
	adder0804: full_adder port map(a => p31(24), b => s696, c_in => p30(25), s => s804, c_out => c804);
	adder0805: full_adder port map(a => c803, b => p28(28), c_in => c804, s => s805, c_out => c805);
	adder0806: full_adder port map(a => p30(26), b => p31(25), c_in => p29(27), s => s806, c_out => c806);
	adder0807: full_adder port map(a => c805, b => p27(30), c_in => c806, s => s807, c_out => c807);
	adder0808: full_adder port map(a => p29(28), b => p30(27), c_in => p28(29), s => s808, c_out => c808);
	adder0809: full_adder port map(a => c807, b => c701, c_in => c808, s => s809, c_out => c809);
	adder0810: full_adder port map(a => p28(30), b => p29(29), c_in => p27(31), s => s810, c_out => c810);
	adder0811: full_adder port map(a => c809, b => p28(31), c_in => c810, s => s811, c_out => c811);
	adder0812: half_adder port map(a => p0(3), b => p1(2), s => s812, c_out => c812);
	adder0813: full_adder port map(a => p2(2), b => p3(1), c_in => c812, s => s813, c_out => c813);
	adder0814: full_adder port map(a => p4(1), b => p5(0), c_in => c813, s => s814, c_out => c814);
	adder0815: full_adder port map(a => p6(0), b => s552, c_in => c814, s => s815, c_out => c815);
	adder0816: full_adder port map(a => s553, b => s554, c_in => c815, s => s816, c_out => c816);
	adder0817: full_adder port map(a => s556, b => s557, c_in => c816, s => s817, c_out => c817);
	adder0818: full_adder port map(a => s559, b => s560, c_in => c817, s => s818, c_out => c818);
	adder0819: full_adder port map(a => s562, b => s563, c_in => c818, s => s819, c_out => c819);
	adder0820: full_adder port map(a => s565, b => s566, c_in => c819, s => s820, c_out => c820);
	adder0821: full_adder port map(a => s568, b => s569, c_in => c820, s => s821, c_out => c821);
	adder0822: full_adder port map(a => s571, b => s572, c_in => c821, s => s822, c_out => c822);
	adder0823: full_adder port map(a => s574, b => s575, c_in => c822, s => s823, c_out => c823);
	adder0824: full_adder port map(a => s577, b => s578, c_in => c823, s => s824, c_out => c824);
	adder0825: full_adder port map(a => s580, b => s581, c_in => c824, s => s825, c_out => c825);
	adder0826: full_adder port map(a => s583, b => s584, c_in => c825, s => s826, c_out => c826);
	adder0827: full_adder port map(a => s586, b => s587, c_in => c826, s => s827, c_out => c827);
	adder0828: full_adder port map(a => s589, b => s590, c_in => c827, s => s828, c_out => c828);
	adder0829: full_adder port map(a => s592, b => s593, c_in => c828, s => s829, c_out => c829);
	adder0830: full_adder port map(a => s595, b => s596, c_in => c829, s => s830, c_out => c830);
	adder0831: full_adder port map(a => s598, b => s599, c_in => c830, s => s831, c_out => c831);
	adder0832: full_adder port map(a => s601, b => s602, c_in => c831, s => s832, c_out => c832);
	adder0833: full_adder port map(a => s604, b => s605, c_in => c832, s => s833, c_out => c833);
	adder0834: full_adder port map(a => s607, b => s608, c_in => c833, s => s834, c_out => c834);
	adder0835: full_adder port map(a => s610, b => s611, c_in => c834, s => s835, c_out => c835);
	adder0836: full_adder port map(a => s613, b => s614, c_in => c835, s => s836, c_out => c836);
	adder0837: full_adder port map(a => s616, b => s617, c_in => c836, s => s837, c_out => c837);
	adder0838: full_adder port map(a => s619, b => s620, c_in => c837, s => s838, c_out => c838);
	adder0839: full_adder port map(a => s622, b => s623, c_in => c838, s => s839, c_out => c839);
	adder0840: full_adder port map(a => s625, b => s626, c_in => c839, s => s840, c_out => c840);
	adder0841: full_adder port map(a => s628, b => s629, c_in => c840, s => s841, c_out => c841);
	adder0842: full_adder port map(a => s631, b => s632, c_in => c841, s => s842, c_out => c842);
	adder0843: full_adder port map(a => s634, b => s635, c_in => c842, s => s843, c_out => c843);
	adder0844: full_adder port map(a => s637, b => s638, c_in => c843, s => s844, c_out => c844);
	adder0845: full_adder port map(a => s640, b => s641, c_in => c844, s => s845, c_out => c845);
	adder0846: full_adder port map(a => s643, b => s644, c_in => c845, s => s846, c_out => c846);
	adder0847: full_adder port map(a => s646, b => s647, c_in => c846, s => s847, c_out => c847);
	adder0848: full_adder port map(a => s649, b => s650, c_in => c847, s => s848, c_out => c848);
	adder0849: full_adder port map(a => s652, b => s653, c_in => c848, s => s849, c_out => c849);
	adder0850: full_adder port map(a => s655, b => s656, c_in => c849, s => s850, c_out => c850);
	adder0851: full_adder port map(a => s658, b => s659, c_in => c850, s => s851, c_out => c851);
	adder0852: full_adder port map(a => s661, b => s662, c_in => c851, s => s852, c_out => c852);
	adder0853: full_adder port map(a => s664, b => s665, c_in => c852, s => s853, c_out => c853);
	adder0854: full_adder port map(a => s667, b => s668, c_in => c853, s => s854, c_out => c854);
	adder0855: full_adder port map(a => s670, b => s671, c_in => c854, s => s855, c_out => c855);
	adder0856: full_adder port map(a => s673, b => s674, c_in => c855, s => s856, c_out => c856);
	adder0857: full_adder port map(a => s676, b => s677, c_in => c856, s => s857, c_out => c857);
	adder0858: full_adder port map(a => s679, b => s680, c_in => c857, s => s858, c_out => c858);
	adder0859: full_adder port map(a => s682, b => s683, c_in => c858, s => s859, c_out => c859);
	adder0860: full_adder port map(a => s685, b => s686, c_in => c859, s => s860, c_out => c860);
	adder0861: full_adder port map(a => s688, b => s689, c_in => c860, s => s861, c_out => c861);
	adder0862: full_adder port map(a => s691, b => s692, c_in => c861, s => s862, c_out => c862);
	adder0863: full_adder port map(a => s694, b => s695, c_in => c862, s => s863, c_out => c863);
	adder0864: full_adder port map(a => s697, b => s698, c_in => c863, s => s864, c_out => c864);
	adder0865: full_adder port map(a => s699, b => s700, c_in => c864, s => s865, c_out => c865);
	adder0866: full_adder port map(a => p31(26), b => s701, c_in => c865, s => s866, c_out => c866);
	adder0867: full_adder port map(a => p30(28), b => p31(27), c_in => c866, s => s867, c_out => c867);
	adder0868: full_adder port map(a => p29(30), b => p30(29), c_in => c867, s => s868, c_out => c868);
	adder0869: full_adder port map(a => c811, b => p29(31), c_in => c868, s => s869, c_out => c869);
	adder0870: half_adder port map(a => p0(2), b => p1(1), s => s870, c_out => c870);
	adder0871: full_adder port map(a => p2(1), b => p3(0), c_in => c870, s => s871, c_out => c871);
	adder0872: full_adder port map(a => p4(0), b => s702, c_in => c871, s => s872, c_out => c872);
	adder0873: full_adder port map(a => s703, b => s704, c_in => c872, s => s873, c_out => c873);
	adder0874: full_adder port map(a => s705, b => s706, c_in => c873, s => s874, c_out => c874);
	adder0875: full_adder port map(a => s707, b => s708, c_in => c874, s => s875, c_out => c875);
	adder0876: full_adder port map(a => s709, b => s710, c_in => c875, s => s876, c_out => c876);
	adder0877: full_adder port map(a => s711, b => s712, c_in => c876, s => s877, c_out => c877);
	adder0878: full_adder port map(a => s713, b => s714, c_in => c877, s => s878, c_out => c878);
	adder0879: full_adder port map(a => s715, b => s716, c_in => c878, s => s879, c_out => c879);
	adder0880: full_adder port map(a => s717, b => s718, c_in => c879, s => s880, c_out => c880);
	adder0881: full_adder port map(a => s719, b => s720, c_in => c880, s => s881, c_out => c881);
	adder0882: full_adder port map(a => s721, b => s722, c_in => c881, s => s882, c_out => c882);
	adder0883: full_adder port map(a => s723, b => s724, c_in => c882, s => s883, c_out => c883);
	adder0884: full_adder port map(a => s725, b => s726, c_in => c883, s => s884, c_out => c884);
	adder0885: full_adder port map(a => s727, b => s728, c_in => c884, s => s885, c_out => c885);
	adder0886: full_adder port map(a => s729, b => s730, c_in => c885, s => s886, c_out => c886);
	adder0887: full_adder port map(a => s731, b => s732, c_in => c886, s => s887, c_out => c887);
	adder0888: full_adder port map(a => s733, b => s734, c_in => c887, s => s888, c_out => c888);
	adder0889: full_adder port map(a => s735, b => s736, c_in => c888, s => s889, c_out => c889);
	adder0890: full_adder port map(a => s737, b => s738, c_in => c889, s => s890, c_out => c890);
	adder0891: full_adder port map(a => s739, b => s740, c_in => c890, s => s891, c_out => c891);
	adder0892: full_adder port map(a => s741, b => s742, c_in => c891, s => s892, c_out => c892);
	adder0893: full_adder port map(a => s743, b => s744, c_in => c892, s => s893, c_out => c893);
	adder0894: full_adder port map(a => s745, b => s746, c_in => c893, s => s894, c_out => c894);
	adder0895: full_adder port map(a => s747, b => s748, c_in => c894, s => s895, c_out => c895);
	adder0896: full_adder port map(a => s749, b => s750, c_in => c895, s => s896, c_out => c896);
	adder0897: full_adder port map(a => s751, b => s752, c_in => c896, s => s897, c_out => c897);
	adder0898: full_adder port map(a => s753, b => s754, c_in => c897, s => s898, c_out => c898);
	adder0899: full_adder port map(a => s755, b => s756, c_in => c898, s => s899, c_out => c899);
	adder0900: full_adder port map(a => s757, b => s758, c_in => c899, s => s900, c_out => c900);
	adder0901: full_adder port map(a => s759, b => s760, c_in => c900, s => s901, c_out => c901);
	adder0902: full_adder port map(a => s761, b => s762, c_in => c901, s => s902, c_out => c902);
	adder0903: full_adder port map(a => s763, b => s764, c_in => c902, s => s903, c_out => c903);
	adder0904: full_adder port map(a => s765, b => s766, c_in => c903, s => s904, c_out => c904);
	adder0905: full_adder port map(a => s767, b => s768, c_in => c904, s => s905, c_out => c905);
	adder0906: full_adder port map(a => s769, b => s770, c_in => c905, s => s906, c_out => c906);
	adder0907: full_adder port map(a => s771, b => s772, c_in => c906, s => s907, c_out => c907);
	adder0908: full_adder port map(a => s773, b => s774, c_in => c907, s => s908, c_out => c908);
	adder0909: full_adder port map(a => s775, b => s776, c_in => c908, s => s909, c_out => c909);
	adder0910: full_adder port map(a => s777, b => s778, c_in => c909, s => s910, c_out => c910);
	adder0911: full_adder port map(a => s779, b => s780, c_in => c910, s => s911, c_out => c911);
	adder0912: full_adder port map(a => s781, b => s782, c_in => c911, s => s912, c_out => c912);
	adder0913: full_adder port map(a => s783, b => s784, c_in => c912, s => s913, c_out => c913);
	adder0914: full_adder port map(a => s785, b => s786, c_in => c913, s => s914, c_out => c914);
	adder0915: full_adder port map(a => s787, b => s788, c_in => c914, s => s915, c_out => c915);
	adder0916: full_adder port map(a => s789, b => s790, c_in => c915, s => s916, c_out => c916);
	adder0917: full_adder port map(a => s791, b => s792, c_in => c916, s => s917, c_out => c917);
	adder0918: full_adder port map(a => s793, b => s794, c_in => c917, s => s918, c_out => c918);
	adder0919: full_adder port map(a => s795, b => s796, c_in => c918, s => s919, c_out => c919);
	adder0920: full_adder port map(a => s797, b => s798, c_in => c919, s => s920, c_out => c920);
	adder0921: full_adder port map(a => s799, b => s800, c_in => c920, s => s921, c_out => c921);
	adder0922: full_adder port map(a => s801, b => s802, c_in => c921, s => s922, c_out => c922);
	adder0923: full_adder port map(a => s803, b => s804, c_in => c922, s => s923, c_out => c923);
	adder0924: full_adder port map(a => s805, b => s806, c_in => c923, s => s924, c_out => c924);
	adder0925: full_adder port map(a => s807, b => s808, c_in => c924, s => s925, c_out => c925);
	adder0926: full_adder port map(a => s809, b => s810, c_in => c925, s => s926, c_out => c926);
	adder0927: full_adder port map(a => p31(28), b => s811, c_in => c926, s => s927, c_out => c927);
	adder0928: full_adder port map(a => p30(30), b => p31(29), c_in => c927, s => s928, c_out => c928);
	adder0929: full_adder port map(a => c869, b => p30(31), c_in => c928, s => s929, c_out => c929);
	flipf0930: flip_flop port map(clk => clk, rst => rst, ce => ce, d => p0(0), q => f0);
	flipf0931: flip_flop port map(clk => clk, rst => rst, ce => ce, d => p0(1), q => f1);
	flipf0932: flip_flop port map(clk => clk, rst => rst, ce => ce, d => p1(0), q => f2);
	flipf0933: flip_flop port map(clk => clk, rst => rst, ce => ce, d => p2(0), q => f3);
	flipf0934: flip_flop port map(clk => clk, rst => rst, ce => ce, d => s870, q => f4);
	flipf0935: flip_flop port map(clk => clk, rst => rst, ce => ce, d => s812, q => f5);
	flipf0936: flip_flop port map(clk => clk, rst => rst, ce => ce, d => s871, q => f6);
	flipf0937: flip_flop port map(clk => clk, rst => rst, ce => ce, d => s813, q => f7);
	flipf0938: flip_flop port map(clk => clk, rst => rst, ce => ce, d => s872, q => f8);
	flipf0939: flip_flop port map(clk => clk, rst => rst, ce => ce, d => s814, q => f9);
	flipf0940: flip_flop port map(clk => clk, rst => rst, ce => ce, d => s873, q => f10);
	flipf0941: flip_flop port map(clk => clk, rst => rst, ce => ce, d => s815, q => f11);
	flipf0942: flip_flop port map(clk => clk, rst => rst, ce => ce, d => s874, q => f12);
	flipf0943: flip_flop port map(clk => clk, rst => rst, ce => ce, d => s816, q => f13);
	flipf0944: flip_flop port map(clk => clk, rst => rst, ce => ce, d => s875, q => f14);
	flipf0945: flip_flop port map(clk => clk, rst => rst, ce => ce, d => s817, q => f15);
	flipf0946: flip_flop port map(clk => clk, rst => rst, ce => ce, d => s876, q => f16);
	flipf0947: flip_flop port map(clk => clk, rst => rst, ce => ce, d => s818, q => f17);
	flipf0948: flip_flop port map(clk => clk, rst => rst, ce => ce, d => s877, q => f18);
	flipf0949: flip_flop port map(clk => clk, rst => rst, ce => ce, d => s819, q => f19);
	flipf0950: flip_flop port map(clk => clk, rst => rst, ce => ce, d => s878, q => f20);
	flipf0951: flip_flop port map(clk => clk, rst => rst, ce => ce, d => s820, q => f21);
	flipf0952: flip_flop port map(clk => clk, rst => rst, ce => ce, d => s879, q => f22);
	flipf0953: flip_flop port map(clk => clk, rst => rst, ce => ce, d => s821, q => f23);
	flipf0954: flip_flop port map(clk => clk, rst => rst, ce => ce, d => s880, q => f24);
	flipf0955: flip_flop port map(clk => clk, rst => rst, ce => ce, d => s822, q => f25);
	flipf0956: flip_flop port map(clk => clk, rst => rst, ce => ce, d => s881, q => f26);
	flipf0957: flip_flop port map(clk => clk, rst => rst, ce => ce, d => s823, q => f27);
	flipf0958: flip_flop port map(clk => clk, rst => rst, ce => ce, d => s882, q => f28);
	flipf0959: flip_flop port map(clk => clk, rst => rst, ce => ce, d => s824, q => f29);
	flipf0960: flip_flop port map(clk => clk, rst => rst, ce => ce, d => s883, q => f30);
	flipf0961: flip_flop port map(clk => clk, rst => rst, ce => ce, d => s825, q => f31);
	flipf0962: flip_flop port map(clk => clk, rst => rst, ce => ce, d => s884, q => f32);
	flipf0963: flip_flop port map(clk => clk, rst => rst, ce => ce, d => s826, q => f33);
	flipf0964: flip_flop port map(clk => clk, rst => rst, ce => ce, d => s885, q => f34);
	flipf0965: flip_flop port map(clk => clk, rst => rst, ce => ce, d => s827, q => f35);
	flipf0966: flip_flop port map(clk => clk, rst => rst, ce => ce, d => s886, q => f36);
	flipf0967: flip_flop port map(clk => clk, rst => rst, ce => ce, d => s828, q => f37);
	flipf0968: flip_flop port map(clk => clk, rst => rst, ce => ce, d => s887, q => f38);
	flipf0969: flip_flop port map(clk => clk, rst => rst, ce => ce, d => s829, q => f39);
	flipf0970: flip_flop port map(clk => clk, rst => rst, ce => ce, d => s888, q => f40);
	flipf0971: flip_flop port map(clk => clk, rst => rst, ce => ce, d => s830, q => f41);
	flipf0972: flip_flop port map(clk => clk, rst => rst, ce => ce, d => s889, q => f42);
	flipf0973: flip_flop port map(clk => clk, rst => rst, ce => ce, d => s831, q => f43);
	flipf0974: flip_flop port map(clk => clk, rst => rst, ce => ce, d => s890, q => f44);
	flipf0975: flip_flop port map(clk => clk, rst => rst, ce => ce, d => s832, q => f45);
	flipf0976: flip_flop port map(clk => clk, rst => rst, ce => ce, d => s891, q => f46);
	flipf0977: flip_flop port map(clk => clk, rst => rst, ce => ce, d => s833, q => f47);
	flipf0978: flip_flop port map(clk => clk, rst => rst, ce => ce, d => s892, q => f48);
	flipf0979: flip_flop port map(clk => clk, rst => rst, ce => ce, d => s834, q => f49);
	flipf0980: flip_flop port map(clk => clk, rst => rst, ce => ce, d => s893, q => f50);
	flipf0981: flip_flop port map(clk => clk, rst => rst, ce => ce, d => s835, q => f51);
	flipf0982: flip_flop port map(clk => clk, rst => rst, ce => ce, d => s894, q => f52);
	flipf0983: flip_flop port map(clk => clk, rst => rst, ce => ce, d => s836, q => f53);
	flipf0984: flip_flop port map(clk => clk, rst => rst, ce => ce, d => s895, q => f54);
	flipf0985: flip_flop port map(clk => clk, rst => rst, ce => ce, d => s837, q => f55);
	flipf0986: flip_flop port map(clk => clk, rst => rst, ce => ce, d => s896, q => f56);
	flipf0987: flip_flop port map(clk => clk, rst => rst, ce => ce, d => s838, q => f57);
	flipf0988: flip_flop port map(clk => clk, rst => rst, ce => ce, d => s897, q => f58);
	flipf0989: flip_flop port map(clk => clk, rst => rst, ce => ce, d => s839, q => f59);
	flipf0990: flip_flop port map(clk => clk, rst => rst, ce => ce, d => s898, q => f60);
	flipf0991: flip_flop port map(clk => clk, rst => rst, ce => ce, d => s840, q => f61);
	flipf0992: flip_flop port map(clk => clk, rst => rst, ce => ce, d => s899, q => f62);
	flipf0993: flip_flop port map(clk => clk, rst => rst, ce => ce, d => s841, q => f63);
	flipf0994: flip_flop port map(clk => clk, rst => rst, ce => ce, d => s900, q => f64);
	flipf0995: flip_flop port map(clk => clk, rst => rst, ce => ce, d => s842, q => f65);
	flipf0996: flip_flop port map(clk => clk, rst => rst, ce => ce, d => s901, q => f66);
	flipf0997: flip_flop port map(clk => clk, rst => rst, ce => ce, d => s843, q => f67);
	flipf0998: flip_flop port map(clk => clk, rst => rst, ce => ce, d => s902, q => f68);
	flipf0999: flip_flop port map(clk => clk, rst => rst, ce => ce, d => s844, q => f69);
	flipf1000: flip_flop port map(clk => clk, rst => rst, ce => ce, d => s903, q => f70);
	flipf1001: flip_flop port map(clk => clk, rst => rst, ce => ce, d => s845, q => f71);
	flipf1002: flip_flop port map(clk => clk, rst => rst, ce => ce, d => s904, q => f72);
	flipf1003: flip_flop port map(clk => clk, rst => rst, ce => ce, d => s846, q => f73);
	flipf1004: flip_flop port map(clk => clk, rst => rst, ce => ce, d => s905, q => f74);
	flipf1005: flip_flop port map(clk => clk, rst => rst, ce => ce, d => s847, q => f75);
	flipf1006: flip_flop port map(clk => clk, rst => rst, ce => ce, d => s906, q => f76);
	flipf1007: flip_flop port map(clk => clk, rst => rst, ce => ce, d => s848, q => f77);
	flipf1008: flip_flop port map(clk => clk, rst => rst, ce => ce, d => s907, q => f78);
	flipf1009: flip_flop port map(clk => clk, rst => rst, ce => ce, d => s849, q => f79);
	flipf1010: flip_flop port map(clk => clk, rst => rst, ce => ce, d => s908, q => f80);
	flipf1011: flip_flop port map(clk => clk, rst => rst, ce => ce, d => s850, q => f81);
	flipf1012: flip_flop port map(clk => clk, rst => rst, ce => ce, d => s909, q => f82);
	flipf1013: flip_flop port map(clk => clk, rst => rst, ce => ce, d => s851, q => f83);
	flipf1014: flip_flop port map(clk => clk, rst => rst, ce => ce, d => s910, q => f84);
	flipf1015: flip_flop port map(clk => clk, rst => rst, ce => ce, d => s852, q => f85);
	flipf1016: flip_flop port map(clk => clk, rst => rst, ce => ce, d => s911, q => f86);
	flipf1017: flip_flop port map(clk => clk, rst => rst, ce => ce, d => s853, q => f87);
	flipf1018: flip_flop port map(clk => clk, rst => rst, ce => ce, d => s912, q => f88);
	flipf1019: flip_flop port map(clk => clk, rst => rst, ce => ce, d => s854, q => f89);
	flipf1020: flip_flop port map(clk => clk, rst => rst, ce => ce, d => s913, q => f90);
	flipf1021: flip_flop port map(clk => clk, rst => rst, ce => ce, d => s855, q => f91);
	flipf1022: flip_flop port map(clk => clk, rst => rst, ce => ce, d => s914, q => f92);
	flipf1023: flip_flop port map(clk => clk, rst => rst, ce => ce, d => s856, q => f93);
	flipf1024: flip_flop port map(clk => clk, rst => rst, ce => ce, d => s915, q => f94);
	flipf1025: flip_flop port map(clk => clk, rst => rst, ce => ce, d => s857, q => f95);
	flipf1026: flip_flop port map(clk => clk, rst => rst, ce => ce, d => s916, q => f96);
	flipf1027: flip_flop port map(clk => clk, rst => rst, ce => ce, d => s858, q => f97);
	flipf1028: flip_flop port map(clk => clk, rst => rst, ce => ce, d => s917, q => f98);
	flipf1029: flip_flop port map(clk => clk, rst => rst, ce => ce, d => s859, q => f99);
	flipf1030: flip_flop port map(clk => clk, rst => rst, ce => ce, d => s918, q => f100);
	flipf1031: flip_flop port map(clk => clk, rst => rst, ce => ce, d => s860, q => f101);
	flipf1032: flip_flop port map(clk => clk, rst => rst, ce => ce, d => s919, q => f102);
	flipf1033: flip_flop port map(clk => clk, rst => rst, ce => ce, d => s861, q => f103);
	flipf1034: flip_flop port map(clk => clk, rst => rst, ce => ce, d => s920, q => f104);
	flipf1035: flip_flop port map(clk => clk, rst => rst, ce => ce, d => s862, q => f105);
	flipf1036: flip_flop port map(clk => clk, rst => rst, ce => ce, d => s921, q => f106);
	flipf1037: flip_flop port map(clk => clk, rst => rst, ce => ce, d => s863, q => f107);
	flipf1038: flip_flop port map(clk => clk, rst => rst, ce => ce, d => s922, q => f108);
	flipf1039: flip_flop port map(clk => clk, rst => rst, ce => ce, d => s864, q => f109);
	flipf1040: flip_flop port map(clk => clk, rst => rst, ce => ce, d => s923, q => f110);
	flipf1041: flip_flop port map(clk => clk, rst => rst, ce => ce, d => s865, q => f111);
	flipf1042: flip_flop port map(clk => clk, rst => rst, ce => ce, d => s924, q => f112);
	flipf1043: flip_flop port map(clk => clk, rst => rst, ce => ce, d => s866, q => f113);
	flipf1044: flip_flop port map(clk => clk, rst => rst, ce => ce, d => s925, q => f114);
	flipf1045: flip_flop port map(clk => clk, rst => rst, ce => ce, d => s867, q => f115);
	flipf1046: flip_flop port map(clk => clk, rst => rst, ce => ce, d => s926, q => f116);
	flipf1047: flip_flop port map(clk => clk, rst => rst, ce => ce, d => s868, q => f117);
	flipf1048: flip_flop port map(clk => clk, rst => rst, ce => ce, d => s927, q => f118);
	flipf1049: flip_flop port map(clk => clk, rst => rst, ce => ce, d => s869, q => f119);
	flipf1050: flip_flop port map(clk => clk, rst => rst, ce => ce, d => s928, q => f120);
	flipf1051: flip_flop port map(clk => clk, rst => rst, ce => ce, d => p31(30), q => f121);
	flipf1052: flip_flop port map(clk => clk, rst => rst, ce => ce, d => s929, q => f122);
	flipf1053: flip_flop port map(clk => clk, rst => rst, ce => ce, d => c929, q => f123);
	flipf1054: flip_flop port map(clk => clk, rst => rst, ce => ce, d => p31(31), q => f124);
	flipf1055: flip_flop port map(clk => clk, rst => rst, ce => ce, d => sgn, q => f125);
	adder1056: half_adder port map(a => f1, b => f2, s => s930, c_out => c930);
	adder1057: full_adder port map(a => f3, b => f4, c_in => c930, s => s931, c_out => c931);
	adder1058: full_adder port map(a => f5, b => f6, c_in => c931, s => s932, c_out => c932);
	adder1059: full_adder port map(a => f7, b => f8, c_in => c932, s => s933, c_out => c933);
	adder1060: full_adder port map(a => f9, b => f10, c_in => c933, s => s934, c_out => c934);
	adder1061: full_adder port map(a => f11, b => f12, c_in => c934, s => s935, c_out => c935);
	adder1062: full_adder port map(a => f13, b => f14, c_in => c935, s => s936, c_out => c936);
	adder1063: full_adder port map(a => f15, b => f16, c_in => c936, s => s937, c_out => c937);
	adder1064: full_adder port map(a => f17, b => f18, c_in => c937, s => s938, c_out => c938);
	adder1065: full_adder port map(a => f19, b => f20, c_in => c938, s => s939, c_out => c939);
	adder1066: full_adder port map(a => f21, b => f22, c_in => c939, s => s940, c_out => c940);
	adder1067: full_adder port map(a => f23, b => f24, c_in => c940, s => s941, c_out => c941);
	adder1068: full_adder port map(a => f25, b => f26, c_in => c941, s => s942, c_out => c942);
	adder1069: full_adder port map(a => f27, b => f28, c_in => c942, s => s943, c_out => c943);
	adder1070: full_adder port map(a => f29, b => f30, c_in => c943, s => s944, c_out => c944);
	adder1071: full_adder port map(a => f31, b => f32, c_in => c944, s => s945, c_out => c945);
	adder1072: full_adder port map(a => f33, b => f34, c_in => c945, s => s946, c_out => c946);
	adder1073: full_adder port map(a => f35, b => f36, c_in => c946, s => s947, c_out => c947);
	adder1074: full_adder port map(a => f37, b => f38, c_in => c947, s => s948, c_out => c948);
	adder1075: full_adder port map(a => f39, b => f40, c_in => c948, s => s949, c_out => c949);
	adder1076: full_adder port map(a => f41, b => f42, c_in => c949, s => s950, c_out => c950);
	adder1077: full_adder port map(a => f43, b => f44, c_in => c950, s => s951, c_out => c951);
	adder1078: full_adder port map(a => f45, b => f46, c_in => c951, s => s952, c_out => c952);
	adder1079: full_adder port map(a => f47, b => f48, c_in => c952, s => s953, c_out => c953);
	adder1080: full_adder port map(a => f49, b => f50, c_in => c953, s => s954, c_out => c954);
	adder1081: full_adder port map(a => f51, b => f52, c_in => c954, s => s955, c_out => c955);
	adder1082: full_adder port map(a => f53, b => f54, c_in => c955, s => s956, c_out => c956);
	adder1083: full_adder port map(a => f55, b => f56, c_in => c956, s => s957, c_out => c957);
	adder1084: full_adder port map(a => f57, b => f58, c_in => c957, s => s958, c_out => c958);
	adder1085: full_adder port map(a => f59, b => f60, c_in => c958, s => s959, c_out => c959);
	adder1086: full_adder port map(a => f61, b => f62, c_in => c959, s => s960, c_out => c960);
	adder1087: full_adder port map(a => f63, b => f64, c_in => c960, s => s961, c_out => c961);
	adder1088: full_adder port map(a => f65, b => f66, c_in => c961, s => s962, c_out => c962);
	adder1089: full_adder port map(a => f67, b => f68, c_in => c962, s => s963, c_out => c963);
	adder1090: full_adder port map(a => f69, b => f70, c_in => c963, s => s964, c_out => c964);
	adder1091: full_adder port map(a => f71, b => f72, c_in => c964, s => s965, c_out => c965);
	adder1092: full_adder port map(a => f73, b => f74, c_in => c965, s => s966, c_out => c966);
	adder1093: full_adder port map(a => f75, b => f76, c_in => c966, s => s967, c_out => c967);
	adder1094: full_adder port map(a => f77, b => f78, c_in => c967, s => s968, c_out => c968);
	adder1095: full_adder port map(a => f79, b => f80, c_in => c968, s => s969, c_out => c969);
	adder1096: full_adder port map(a => f81, b => f82, c_in => c969, s => s970, c_out => c970);
	adder1097: full_adder port map(a => f83, b => f84, c_in => c970, s => s971, c_out => c971);
	adder1098: full_adder port map(a => f85, b => f86, c_in => c971, s => s972, c_out => c972);
	adder1099: full_adder port map(a => f87, b => f88, c_in => c972, s => s973, c_out => c973);
	adder1100: full_adder port map(a => f89, b => f90, c_in => c973, s => s974, c_out => c974);
	adder1101: full_adder port map(a => f91, b => f92, c_in => c974, s => s975, c_out => c975);
	adder1102: full_adder port map(a => f93, b => f94, c_in => c975, s => s976, c_out => c976);
	adder1103: full_adder port map(a => f95, b => f96, c_in => c976, s => s977, c_out => c977);
	adder1104: full_adder port map(a => f97, b => f98, c_in => c977, s => s978, c_out => c978);
	adder1105: full_adder port map(a => f99, b => f100, c_in => c978, s => s979, c_out => c979);
	adder1106: full_adder port map(a => f101, b => f102, c_in => c979, s => s980, c_out => c980);
	adder1107: full_adder port map(a => f103, b => f104, c_in => c980, s => s981, c_out => c981);
	adder1108: full_adder port map(a => f105, b => f106, c_in => c981, s => s982, c_out => c982);
	adder1109: full_adder port map(a => f107, b => f108, c_in => c982, s => s983, c_out => c983);
	adder1110: full_adder port map(a => f109, b => f110, c_in => c983, s => s984, c_out => c984);
	adder1111: full_adder port map(a => f111, b => f112, c_in => c984, s => s985, c_out => c985);
	adder1112: full_adder port map(a => f113, b => f114, c_in => c985, s => s986, c_out => c986);
	adder1113: full_adder port map(a => f115, b => f116, c_in => c986, s => s987, c_out => c987);
	adder1114: full_adder port map(a => f117, b => f118, c_in => c987, s => s988, c_out => c988);
	adder1115: full_adder port map(a => f119, b => f120, c_in => c988, s => s989, c_out => c989);
	adder1116: full_adder port map(a => f121, b => f122, c_in => c989, s => s990, c_out => c990);
	adder1117: full_adder port map(a => f123, b => f124, c_in => c990, s => s991, c_out => c991);
	adder1118: half_adder port map(a => c991, b => f125, s => s992, c_out => c992);

	c_mult <= s992 & s991 & s990 & s989 & s988 & s987 & s986 & s985 & s984 & s983 & s982 & s981 & s980 & s979 & s978 & s977 & s976 & s975 & s974 & s973 & s972 & s971 & s970 & s969 & s968 & s967 & s966 & s965 & s964 & s963 & s962 & s961 & s960 & s959 & s958 & s957 & s956 & s955 & s954 & s953 & s952 & s951 & s950 & s949 & s948 & s947 & s946 & s945 & s944 & s943 & s942 & s941 & s940 & s939 & s938 & s937 & s936 & s935 & s934 & s933 & s932 & s931 & s930 & f0;
end;
